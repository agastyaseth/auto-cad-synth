// `include "adder32.v"
// `include "mult32.v"
module PE (input [31:0] x, input [31:0] w, input [31:0] acc, output reg [31:0] res, input clk, output reg [31:0] wout);
  
  reg [31:0] S1;
  
  wire [31:0] addout,multout;
  always @(posedge clk) begin
    res <= addout;
   // res <= S1;
    wout <= w;
  end
  
mult32 m1(.clk(clk),.en(1'b1),.rst(1'b0),.a(x),.b(w),.z(multout),.output_ready());
adder32 a1(.clk(clk),.en(1'b1),.rst(1'b0),.a(multout),.b(acc),.z(addout),.output_ready());
endmodule

module systolicfull_128(input [31:0] x0,input [31:0] x1,input [31:0] x2,input [31:0] x3,input [31:0] x4,input [31:0] x5,input [31:0] x6,input [31:0] x7,input [31:0] x8,input [31:0] x9,input [31:0] x10,input [31:0] x11,input [31:0] x12,input [31:0] x13,input [31:0] x14,input [31:0] x15,input [31:0] x16,
	input [31:0] x17,input [31:0] x18,input [31:0] x19,input [31:0] x20,input [31:0] x21,input [31:0] x22,input [31:0] x23,input [31:0] x24,input [31:0] x25,input [31:0] x26,input [31:0] x27,input [31:0] x28,input [31:0] x29,input [31:0] x30,input [31:0] x31,input [31:0] x32,
	input [31:0] x33,input [31:0] x34,input [31:0] x35,input [31:0] x36,input [31:0] x37,input [31:0] x38,input [31:0] x39,input [31:0] x40,input [31:0] x41,input [31:0] x42,input [31:0] x43,input [31:0] x44,input [31:0] x45,input [31:0] x46,input [31:0] x47,input [31:0] x48,
	input [31:0] x49,input [31:0] x50,input [31:0] x51,input [31:0] x52,input [31:0] x53,input [31:0] x54,input [31:0] x55,input [31:0] x56,input [31:0] x57,input [31:0] x58,input [31:0] x59,input [31:0] x60,input [31:0] x61,input [31:0] x62,input [31:0] x63,input [31:0] x64,
	input [31:0] x65,input [31:0] x66,input [31:0] x67,input [31:0] x68,input [31:0] x69,input [31:0] x70,input [31:0] x71,input [31:0] x72,input [31:0] x73,input [31:0] x74,input [31:0] x75,input [31:0] x76,input [31:0] x77,input [31:0] x78,input [31:0] x79,input [31:0] x80,
	input [31:0] x81,input [31:0] x82,input [31:0] x83,input [31:0] x84,input [31:0] x85,input [31:0] x86,input [31:0] x87,input [31:0] x88,input [31:0] x89,input [31:0] x90,input [31:0] x91,input [31:0] x92,input [31:0] x93,input [31:0] x94,input [31:0] x95,input [31:0] x96,
	input [31:0] x97,input [31:0] x98,input [31:0] x99,input [31:0] x100,input [31:0] x101,input [31:0] x102,input [31:0] x103,input [31:0] x104,input [31:0] x105,input [31:0] x106,input [31:0] x107,input [31:0] x108,input [31:0] x109,input [31:0] x110,input [31:0] x111,input [31:0] x112,
	input [31:0] x113,input [31:0] x114,input [31:0] x115,input [31:0] x116,input [31:0] x117,input [31:0] x118,input [31:0] x119,input [31:0] x120,input [31:0] x121,input [31:0] x122,input [31:0] x123,input [31:0] x124,input [31:0] x125,input [31:0] x126,input [31:0] x127,
	input [31:0] w0,input [31:0] w1,input [31:0] w2,input [31:0] w3,input [31:0] w4,input [31:0] w5,input [31:0] w6,input [31:0] w7,input [31:0] w8,input [31:0] w9,input [31:0] w10,input [31:0] w11,input [31:0] w12,input [31:0] w13,input [31:0] w14,input [31:0] w15,input [31:0] w16,
	input [31:0] w17,input [31:0] w18,input [31:0] w19,input [31:0] w20,input [31:0] w21,input [31:0] w22,input [31:0] w23,input [31:0] w24,input [31:0] w25,input [31:0] w26,input [31:0] w27,input [31:0] w28,input [31:0] w29,input [31:0] w30,input [31:0] w31,input [31:0] w32,
	input [31:0] w33,input [31:0] w34,input [31:0] w35,input [31:0] w36,input [31:0] w37,input [31:0] w38,input [31:0] w39,input [31:0] w40,input [31:0] w41,input [31:0] w42,input [31:0] w43,input [31:0] w44,input [31:0] w45,input [31:0] w46,input [31:0] w47,input [31:0] w48,
	input [31:0] w49,input [31:0] w50,input [31:0] w51,input [31:0] w52,input [31:0] w53,input [31:0] w54,input [31:0] w55,input [31:0] w56,input [31:0] w57,input [31:0] w58,input [31:0] w59,input [31:0] w60,input [31:0] w61,input [31:0] w62,input [31:0] w63,input [31:0] w64,
	input [31:0] w65,input [31:0] w66,input [31:0] w67,input [31:0] w68,input [31:0] w69,input [31:0] w70,input [31:0] w71,input [31:0] w72,input [31:0] w73,input [31:0] w74,input [31:0] w75,input [31:0] w76,input [31:0] w77,input [31:0] w78,input [31:0] w79,input [31:0] w80,
	input [31:0] w81,input [31:0] w82,input [31:0] w83,input [31:0] w84,input [31:0] w85,input [31:0] w86,input [31:0] w87,input [31:0] w88,input [31:0] w89,input [31:0] w90,input [31:0] w91,input [31:0] w92,input [31:0] w93,input [31:0] w94,input [31:0] w95,input [31:0] w96,
	input [31:0] w97,input [31:0] w98,input [31:0] w99,input [31:0] w100,input [31:0] w101,input [31:0] w102,input [31:0] w103,input [31:0] w104,input [31:0] w105,input [31:0] w106,input [31:0] w107,input [31:0] w108,input [31:0] w109,input [31:0] w110,input [31:0] w111,input [31:0] w112,
	input [31:0] w113,input [31:0] w114,input [31:0] w115,input [31:0] w116,input [31:0] w117,input [31:0] w118,input [31:0] w119,input [31:0] w120,input [31:0] w121,input [31:0] w122,input [31:0] w123,input [31:0] w124,input [31:0] w125,input [31:0] w126,input [31:0] w127,
	output [31:0] result0,output [31:0] result1,output [31:0] result2,output [31:0] result3,output [31:0] result4,output [31:0] result5,output [31:0] result6,output [31:0] result7,output [31:0] result8,output [31:0] result9,output [31:0] result10,output [31:0] result11,output [31:0] result12,output [31:0] result13,output [31:0] result14,output [31:0] result15,output [31:0] result16,
	output [31:0] result17,output [31:0] result18,output [31:0] result19,output [31:0] result20,output [31:0] result21,output [31:0] result22,output [31:0] result23,output [31:0] result24,output [31:0] result25,output [31:0] result26,output [31:0] result27,output [31:0] result28,output [31:0] result29,output [31:0] result30,output [31:0] result31,output [31:0] result32,
	output [31:0] result33,output [31:0] result34,output [31:0] result35,output [31:0] result36,output [31:0] result37,output [31:0] result38,output [31:0] result39,output [31:0] result40,output [31:0] result41,output [31:0] result42,output [31:0] result43,output [31:0] result44,output [31:0] result45,output [31:0] result46,output [31:0] result47,output [31:0] result48,
	output [31:0] result49,output [31:0] result50,output [31:0] result51,output [31:0] result52,output [31:0] result53,output [31:0] result54,output [31:0] result55,output [31:0] result56,output [31:0] result57,output [31:0] result58,output [31:0] result59,output [31:0] result60,output [31:0] result61,output [31:0] result62,output [31:0] result63,output [31:0] result64,
	output [31:0] result65,output [31:0] result66,output [31:0] result67,output [31:0] result68,output [31:0] result69,output [31:0] result70,output [31:0] result71,output [31:0] result72,output [31:0] result73,output [31:0] result74,output [31:0] result75,output [31:0] result76,output [31:0] result77,output [31:0] result78,output [31:0] result79,output [31:0] result80,
	output [31:0] result81,output [31:0] result82,output [31:0] result83,output [31:0] result84,output [31:0] result85,output [31:0] result86,output [31:0] result87,output [31:0] result88,output [31:0] result89,output [31:0] result90,output [31:0] result91,output [31:0] result92,output [31:0] result93,output [31:0] result94,output [31:0] result95,output [31:0] result96,
	output [31:0] result97,output [31:0] result98,output [31:0] result99,output [31:0] result100,output [31:0] result101,output [31:0] result102,output [31:0] result103,output [31:0] result104,output [31:0] result105,output [31:0] result106,output [31:0] result107,output [31:0] result108,output [31:0] result109,output [31:0] result110,output [31:0] result111,output [31:0] result112,
	output [31:0] result113,output [31:0] result114,output [31:0] result115,output [31:0] result116,output [31:0] result117,output [31:0] result118,output [31:0] result119,output [31:0] result120,output [31:0] result121,output [31:0] result122,output [31:0] result123,output [31:0] result124,output [31:0] result125,output [31:0] result126,output [31:0] result127,
	output [31:0] weight0,output [31:0] weight1,output [31:0] weight2,output [31:0] weight3,output [31:0] weight4,output [31:0] weight5,output [31:0] weight6,output [31:0] weight7,output [31:0] weight8,output [31:0] weight9,output [31:0] weight10,output [31:0] weight11,output [31:0] weight12,output [31:0] weight13,output [31:0] weight14,output [31:0] weight15,output [31:0] weight16,
	output [31:0] weight17,output [31:0] weight18,output [31:0] weight19,output [31:0] weight20,output [31:0] weight21,output [31:0] weight22,output [31:0] weight23,output [31:0] weight24,output [31:0] weight25,output [31:0] weight26,output [31:0] weight27,output [31:0] weight28,output [31:0] weight29,output [31:0] weight30,output [31:0] weight31,output [31:0] weight32,
	output [31:0] weight33,output [31:0] weight34,output [31:0] weight35,output [31:0] weight36,output [31:0] weight37,output [31:0] weight38,output [31:0] weight39,output [31:0] weight40,output [31:0] weight41,output [31:0] weight42,output [31:0] weight43,output [31:0] weight44,output [31:0] weight45,output [31:0] weight46,output [31:0] weight47,output [31:0] weight48,
	output [31:0] weight49,output [31:0] weight50,output [31:0] weight51,output [31:0] weight52,output [31:0] weight53,output [31:0] weight54,output [31:0] weight55,output [31:0] weight56,output [31:0] weight57,output [31:0] weight58,output [31:0] weight59,output [31:0] weight60,output [31:0] weight61,output [31:0] weight62,output [31:0] weight63,output [31:0] weight64,
	output [31:0] weight65,output [31:0] weight66,output [31:0] weight67,output [31:0] weight68,output [31:0] weight69,output [31:0] weight70,output [31:0] weight71,output [31:0] weight72,output [31:0] weight73,output [31:0] weight74,output [31:0] weight75,output [31:0] weight76,output [31:0] weight77,output [31:0] weight78,output [31:0] weight79,output [31:0] weight80,
	output [31:0] weight81,output [31:0] weight82,output [31:0] weight83,output [31:0] weight84,output [31:0] weight85,output [31:0] weight86,output [31:0] weight87,output [31:0] weight88,output [31:0] weight89,output [31:0] weight90,output [31:0] weight91,output [31:0] weight92,output [31:0] weight93,output [31:0] weight94,output [31:0] weight95,output [31:0] weight96,
	output [31:0] weight97,output [31:0] weight98,output [31:0] weight99,output [31:0] weight100,output [31:0] weight101,output [31:0] weight102,output [31:0] weight103,output [31:0] weight104,output [31:0] weight105,output [31:0] weight106,output [31:0] weight107,output [31:0] weight108,output [31:0] weight109,output [31:0] weight110,output [31:0] weight111,output [31:0] weight112,
	output [31:0] weight113,output [31:0] weight114,output [31:0] weight115,output [31:0] weight116,output [31:0] weight117,output [31:0] weight118,output [31:0] weight119,output [31:0] weight120,output [31:0] weight121,output [31:0] weight122,output [31:0] weight123,output [31:0] weight124,output [31:0] weight125,output [31:0] weight126,output [31:0] weight127,
	input clk); 

	wire [31:0] w0_0,w0_1,w0_2,w0_3,w0_4,w0_5,w0_6,w0_7,w0_8,w0_9,w0_10,w0_11,w0_12,w0_13,w0_14,w0_15,w0_16,
		w0_17,w0_18,w0_19,w0_20,w0_21,w0_22,w0_23,w0_24,w0_25,w0_26,w0_27,w0_28,w0_29,w0_30,w0_31,w0_32,
		w0_33,w0_34,w0_35,w0_36,w0_37,w0_38,w0_39,w0_40,w0_41,w0_42,w0_43,w0_44,w0_45,w0_46,w0_47,w0_48,
		w0_49,w0_50,w0_51,w0_52,w0_53,w0_54,w0_55,w0_56,w0_57,w0_58,w0_59,w0_60,w0_61,w0_62,w0_63,w0_64,
		w0_65,w0_66,w0_67,w0_68,w0_69,w0_70,w0_71,w0_72,w0_73,w0_74,w0_75,w0_76,w0_77,w0_78,w0_79,w0_80,
		w0_81,w0_82,w0_83,w0_84,w0_85,w0_86,w0_87,w0_88,w0_89,w0_90,w0_91,w0_92,w0_93,w0_94,w0_95,w0_96,
		w0_97,w0_98,w0_99,w0_100,w0_101,w0_102,w0_103,w0_104,w0_105,w0_106,w0_107,w0_108,w0_109,w0_110,w0_111,w0_112,
		w0_113,w0_114,w0_115,w0_116,w0_117,w0_118,w0_119,w0_120,w0_121,w0_122,w0_123,w0_124,w0_125,w0_126,
	w1_0,w1_1,w1_2,w1_3,w1_4,w1_5,w1_6,w1_7,w1_8,w1_9,w1_10,w1_11,w1_12,w1_13,w1_14,w1_15,w1_16,
		w1_17,w1_18,w1_19,w1_20,w1_21,w1_22,w1_23,w1_24,w1_25,w1_26,w1_27,w1_28,w1_29,w1_30,w1_31,w1_32,
		w1_33,w1_34,w1_35,w1_36,w1_37,w1_38,w1_39,w1_40,w1_41,w1_42,w1_43,w1_44,w1_45,w1_46,w1_47,w1_48,
		w1_49,w1_50,w1_51,w1_52,w1_53,w1_54,w1_55,w1_56,w1_57,w1_58,w1_59,w1_60,w1_61,w1_62,w1_63,w1_64,
		w1_65,w1_66,w1_67,w1_68,w1_69,w1_70,w1_71,w1_72,w1_73,w1_74,w1_75,w1_76,w1_77,w1_78,w1_79,w1_80,
		w1_81,w1_82,w1_83,w1_84,w1_85,w1_86,w1_87,w1_88,w1_89,w1_90,w1_91,w1_92,w1_93,w1_94,w1_95,w1_96,
		w1_97,w1_98,w1_99,w1_100,w1_101,w1_102,w1_103,w1_104,w1_105,w1_106,w1_107,w1_108,w1_109,w1_110,w1_111,w1_112,
		w1_113,w1_114,w1_115,w1_116,w1_117,w1_118,w1_119,w1_120,w1_121,w1_122,w1_123,w1_124,w1_125,w1_126,
	w2_0,w2_1,w2_2,w2_3,w2_4,w2_5,w2_6,w2_7,w2_8,w2_9,w2_10,w2_11,w2_12,w2_13,w2_14,w2_15,w2_16,
		w2_17,w2_18,w2_19,w2_20,w2_21,w2_22,w2_23,w2_24,w2_25,w2_26,w2_27,w2_28,w2_29,w2_30,w2_31,w2_32,
		w2_33,w2_34,w2_35,w2_36,w2_37,w2_38,w2_39,w2_40,w2_41,w2_42,w2_43,w2_44,w2_45,w2_46,w2_47,w2_48,
		w2_49,w2_50,w2_51,w2_52,w2_53,w2_54,w2_55,w2_56,w2_57,w2_58,w2_59,w2_60,w2_61,w2_62,w2_63,w2_64,
		w2_65,w2_66,w2_67,w2_68,w2_69,w2_70,w2_71,w2_72,w2_73,w2_74,w2_75,w2_76,w2_77,w2_78,w2_79,w2_80,
		w2_81,w2_82,w2_83,w2_84,w2_85,w2_86,w2_87,w2_88,w2_89,w2_90,w2_91,w2_92,w2_93,w2_94,w2_95,w2_96,
		w2_97,w2_98,w2_99,w2_100,w2_101,w2_102,w2_103,w2_104,w2_105,w2_106,w2_107,w2_108,w2_109,w2_110,w2_111,w2_112,
		w2_113,w2_114,w2_115,w2_116,w2_117,w2_118,w2_119,w2_120,w2_121,w2_122,w2_123,w2_124,w2_125,w2_126,
	w3_0,w3_1,w3_2,w3_3,w3_4,w3_5,w3_6,w3_7,w3_8,w3_9,w3_10,w3_11,w3_12,w3_13,w3_14,w3_15,w3_16,
		w3_17,w3_18,w3_19,w3_20,w3_21,w3_22,w3_23,w3_24,w3_25,w3_26,w3_27,w3_28,w3_29,w3_30,w3_31,w3_32,
		w3_33,w3_34,w3_35,w3_36,w3_37,w3_38,w3_39,w3_40,w3_41,w3_42,w3_43,w3_44,w3_45,w3_46,w3_47,w3_48,
		w3_49,w3_50,w3_51,w3_52,w3_53,w3_54,w3_55,w3_56,w3_57,w3_58,w3_59,w3_60,w3_61,w3_62,w3_63,w3_64,
		w3_65,w3_66,w3_67,w3_68,w3_69,w3_70,w3_71,w3_72,w3_73,w3_74,w3_75,w3_76,w3_77,w3_78,w3_79,w3_80,
		w3_81,w3_82,w3_83,w3_84,w3_85,w3_86,w3_87,w3_88,w3_89,w3_90,w3_91,w3_92,w3_93,w3_94,w3_95,w3_96,
		w3_97,w3_98,w3_99,w3_100,w3_101,w3_102,w3_103,w3_104,w3_105,w3_106,w3_107,w3_108,w3_109,w3_110,w3_111,w3_112,
		w3_113,w3_114,w3_115,w3_116,w3_117,w3_118,w3_119,w3_120,w3_121,w3_122,w3_123,w3_124,w3_125,w3_126,
	w4_0,w4_1,w4_2,w4_3,w4_4,w4_5,w4_6,w4_7,w4_8,w4_9,w4_10,w4_11,w4_12,w4_13,w4_14,w4_15,w4_16,
		w4_17,w4_18,w4_19,w4_20,w4_21,w4_22,w4_23,w4_24,w4_25,w4_26,w4_27,w4_28,w4_29,w4_30,w4_31,w4_32,
		w4_33,w4_34,w4_35,w4_36,w4_37,w4_38,w4_39,w4_40,w4_41,w4_42,w4_43,w4_44,w4_45,w4_46,w4_47,w4_48,
		w4_49,w4_50,w4_51,w4_52,w4_53,w4_54,w4_55,w4_56,w4_57,w4_58,w4_59,w4_60,w4_61,w4_62,w4_63,w4_64,
		w4_65,w4_66,w4_67,w4_68,w4_69,w4_70,w4_71,w4_72,w4_73,w4_74,w4_75,w4_76,w4_77,w4_78,w4_79,w4_80,
		w4_81,w4_82,w4_83,w4_84,w4_85,w4_86,w4_87,w4_88,w4_89,w4_90,w4_91,w4_92,w4_93,w4_94,w4_95,w4_96,
		w4_97,w4_98,w4_99,w4_100,w4_101,w4_102,w4_103,w4_104,w4_105,w4_106,w4_107,w4_108,w4_109,w4_110,w4_111,w4_112,
		w4_113,w4_114,w4_115,w4_116,w4_117,w4_118,w4_119,w4_120,w4_121,w4_122,w4_123,w4_124,w4_125,w4_126,
	w5_0,w5_1,w5_2,w5_3,w5_4,w5_5,w5_6,w5_7,w5_8,w5_9,w5_10,w5_11,w5_12,w5_13,w5_14,w5_15,w5_16,
		w5_17,w5_18,w5_19,w5_20,w5_21,w5_22,w5_23,w5_24,w5_25,w5_26,w5_27,w5_28,w5_29,w5_30,w5_31,w5_32,
		w5_33,w5_34,w5_35,w5_36,w5_37,w5_38,w5_39,w5_40,w5_41,w5_42,w5_43,w5_44,w5_45,w5_46,w5_47,w5_48,
		w5_49,w5_50,w5_51,w5_52,w5_53,w5_54,w5_55,w5_56,w5_57,w5_58,w5_59,w5_60,w5_61,w5_62,w5_63,w5_64,
		w5_65,w5_66,w5_67,w5_68,w5_69,w5_70,w5_71,w5_72,w5_73,w5_74,w5_75,w5_76,w5_77,w5_78,w5_79,w5_80,
		w5_81,w5_82,w5_83,w5_84,w5_85,w5_86,w5_87,w5_88,w5_89,w5_90,w5_91,w5_92,w5_93,w5_94,w5_95,w5_96,
		w5_97,w5_98,w5_99,w5_100,w5_101,w5_102,w5_103,w5_104,w5_105,w5_106,w5_107,w5_108,w5_109,w5_110,w5_111,w5_112,
		w5_113,w5_114,w5_115,w5_116,w5_117,w5_118,w5_119,w5_120,w5_121,w5_122,w5_123,w5_124,w5_125,w5_126,
	w6_0,w6_1,w6_2,w6_3,w6_4,w6_5,w6_6,w6_7,w6_8,w6_9,w6_10,w6_11,w6_12,w6_13,w6_14,w6_15,w6_16,
		w6_17,w6_18,w6_19,w6_20,w6_21,w6_22,w6_23,w6_24,w6_25,w6_26,w6_27,w6_28,w6_29,w6_30,w6_31,w6_32,
		w6_33,w6_34,w6_35,w6_36,w6_37,w6_38,w6_39,w6_40,w6_41,w6_42,w6_43,w6_44,w6_45,w6_46,w6_47,w6_48,
		w6_49,w6_50,w6_51,w6_52,w6_53,w6_54,w6_55,w6_56,w6_57,w6_58,w6_59,w6_60,w6_61,w6_62,w6_63,w6_64,
		w6_65,w6_66,w6_67,w6_68,w6_69,w6_70,w6_71,w6_72,w6_73,w6_74,w6_75,w6_76,w6_77,w6_78,w6_79,w6_80,
		w6_81,w6_82,w6_83,w6_84,w6_85,w6_86,w6_87,w6_88,w6_89,w6_90,w6_91,w6_92,w6_93,w6_94,w6_95,w6_96,
		w6_97,w6_98,w6_99,w6_100,w6_101,w6_102,w6_103,w6_104,w6_105,w6_106,w6_107,w6_108,w6_109,w6_110,w6_111,w6_112,
		w6_113,w6_114,w6_115,w6_116,w6_117,w6_118,w6_119,w6_120,w6_121,w6_122,w6_123,w6_124,w6_125,w6_126,
	w7_0,w7_1,w7_2,w7_3,w7_4,w7_5,w7_6,w7_7,w7_8,w7_9,w7_10,w7_11,w7_12,w7_13,w7_14,w7_15,w7_16,
		w7_17,w7_18,w7_19,w7_20,w7_21,w7_22,w7_23,w7_24,w7_25,w7_26,w7_27,w7_28,w7_29,w7_30,w7_31,w7_32,
		w7_33,w7_34,w7_35,w7_36,w7_37,w7_38,w7_39,w7_40,w7_41,w7_42,w7_43,w7_44,w7_45,w7_46,w7_47,w7_48,
		w7_49,w7_50,w7_51,w7_52,w7_53,w7_54,w7_55,w7_56,w7_57,w7_58,w7_59,w7_60,w7_61,w7_62,w7_63,w7_64,
		w7_65,w7_66,w7_67,w7_68,w7_69,w7_70,w7_71,w7_72,w7_73,w7_74,w7_75,w7_76,w7_77,w7_78,w7_79,w7_80,
		w7_81,w7_82,w7_83,w7_84,w7_85,w7_86,w7_87,w7_88,w7_89,w7_90,w7_91,w7_92,w7_93,w7_94,w7_95,w7_96,
		w7_97,w7_98,w7_99,w7_100,w7_101,w7_102,w7_103,w7_104,w7_105,w7_106,w7_107,w7_108,w7_109,w7_110,w7_111,w7_112,
		w7_113,w7_114,w7_115,w7_116,w7_117,w7_118,w7_119,w7_120,w7_121,w7_122,w7_123,w7_124,w7_125,w7_126,
	w8_0,w8_1,w8_2,w8_3,w8_4,w8_5,w8_6,w8_7,w8_8,w8_9,w8_10,w8_11,w8_12,w8_13,w8_14,w8_15,w8_16,
		w8_17,w8_18,w8_19,w8_20,w8_21,w8_22,w8_23,w8_24,w8_25,w8_26,w8_27,w8_28,w8_29,w8_30,w8_31,w8_32,
		w8_33,w8_34,w8_35,w8_36,w8_37,w8_38,w8_39,w8_40,w8_41,w8_42,w8_43,w8_44,w8_45,w8_46,w8_47,w8_48,
		w8_49,w8_50,w8_51,w8_52,w8_53,w8_54,w8_55,w8_56,w8_57,w8_58,w8_59,w8_60,w8_61,w8_62,w8_63,w8_64,
		w8_65,w8_66,w8_67,w8_68,w8_69,w8_70,w8_71,w8_72,w8_73,w8_74,w8_75,w8_76,w8_77,w8_78,w8_79,w8_80,
		w8_81,w8_82,w8_83,w8_84,w8_85,w8_86,w8_87,w8_88,w8_89,w8_90,w8_91,w8_92,w8_93,w8_94,w8_95,w8_96,
		w8_97,w8_98,w8_99,w8_100,w8_101,w8_102,w8_103,w8_104,w8_105,w8_106,w8_107,w8_108,w8_109,w8_110,w8_111,w8_112,
		w8_113,w8_114,w8_115,w8_116,w8_117,w8_118,w8_119,w8_120,w8_121,w8_122,w8_123,w8_124,w8_125,w8_126,
	w9_0,w9_1,w9_2,w9_3,w9_4,w9_5,w9_6,w9_7,w9_8,w9_9,w9_10,w9_11,w9_12,w9_13,w9_14,w9_15,w9_16,
		w9_17,w9_18,w9_19,w9_20,w9_21,w9_22,w9_23,w9_24,w9_25,w9_26,w9_27,w9_28,w9_29,w9_30,w9_31,w9_32,
		w9_33,w9_34,w9_35,w9_36,w9_37,w9_38,w9_39,w9_40,w9_41,w9_42,w9_43,w9_44,w9_45,w9_46,w9_47,w9_48,
		w9_49,w9_50,w9_51,w9_52,w9_53,w9_54,w9_55,w9_56,w9_57,w9_58,w9_59,w9_60,w9_61,w9_62,w9_63,w9_64,
		w9_65,w9_66,w9_67,w9_68,w9_69,w9_70,w9_71,w9_72,w9_73,w9_74,w9_75,w9_76,w9_77,w9_78,w9_79,w9_80,
		w9_81,w9_82,w9_83,w9_84,w9_85,w9_86,w9_87,w9_88,w9_89,w9_90,w9_91,w9_92,w9_93,w9_94,w9_95,w9_96,
		w9_97,w9_98,w9_99,w9_100,w9_101,w9_102,w9_103,w9_104,w9_105,w9_106,w9_107,w9_108,w9_109,w9_110,w9_111,w9_112,
		w9_113,w9_114,w9_115,w9_116,w9_117,w9_118,w9_119,w9_120,w9_121,w9_122,w9_123,w9_124,w9_125,w9_126,
	w10_0,w10_1,w10_2,w10_3,w10_4,w10_5,w10_6,w10_7,w10_8,w10_9,w10_10,w10_11,w10_12,w10_13,w10_14,w10_15,w10_16,
		w10_17,w10_18,w10_19,w10_20,w10_21,w10_22,w10_23,w10_24,w10_25,w10_26,w10_27,w10_28,w10_29,w10_30,w10_31,w10_32,
		w10_33,w10_34,w10_35,w10_36,w10_37,w10_38,w10_39,w10_40,w10_41,w10_42,w10_43,w10_44,w10_45,w10_46,w10_47,w10_48,
		w10_49,w10_50,w10_51,w10_52,w10_53,w10_54,w10_55,w10_56,w10_57,w10_58,w10_59,w10_60,w10_61,w10_62,w10_63,w10_64,
		w10_65,w10_66,w10_67,w10_68,w10_69,w10_70,w10_71,w10_72,w10_73,w10_74,w10_75,w10_76,w10_77,w10_78,w10_79,w10_80,
		w10_81,w10_82,w10_83,w10_84,w10_85,w10_86,w10_87,w10_88,w10_89,w10_90,w10_91,w10_92,w10_93,w10_94,w10_95,w10_96,
		w10_97,w10_98,w10_99,w10_100,w10_101,w10_102,w10_103,w10_104,w10_105,w10_106,w10_107,w10_108,w10_109,w10_110,w10_111,w10_112,
		w10_113,w10_114,w10_115,w10_116,w10_117,w10_118,w10_119,w10_120,w10_121,w10_122,w10_123,w10_124,w10_125,w10_126,
	w11_0,w11_1,w11_2,w11_3,w11_4,w11_5,w11_6,w11_7,w11_8,w11_9,w11_10,w11_11,w11_12,w11_13,w11_14,w11_15,w11_16,
		w11_17,w11_18,w11_19,w11_20,w11_21,w11_22,w11_23,w11_24,w11_25,w11_26,w11_27,w11_28,w11_29,w11_30,w11_31,w11_32,
		w11_33,w11_34,w11_35,w11_36,w11_37,w11_38,w11_39,w11_40,w11_41,w11_42,w11_43,w11_44,w11_45,w11_46,w11_47,w11_48,
		w11_49,w11_50,w11_51,w11_52,w11_53,w11_54,w11_55,w11_56,w11_57,w11_58,w11_59,w11_60,w11_61,w11_62,w11_63,w11_64,
		w11_65,w11_66,w11_67,w11_68,w11_69,w11_70,w11_71,w11_72,w11_73,w11_74,w11_75,w11_76,w11_77,w11_78,w11_79,w11_80,
		w11_81,w11_82,w11_83,w11_84,w11_85,w11_86,w11_87,w11_88,w11_89,w11_90,w11_91,w11_92,w11_93,w11_94,w11_95,w11_96,
		w11_97,w11_98,w11_99,w11_100,w11_101,w11_102,w11_103,w11_104,w11_105,w11_106,w11_107,w11_108,w11_109,w11_110,w11_111,w11_112,
		w11_113,w11_114,w11_115,w11_116,w11_117,w11_118,w11_119,w11_120,w11_121,w11_122,w11_123,w11_124,w11_125,w11_126,
	w12_0,w12_1,w12_2,w12_3,w12_4,w12_5,w12_6,w12_7,w12_8,w12_9,w12_10,w12_11,w12_12,w12_13,w12_14,w12_15,w12_16,
		w12_17,w12_18,w12_19,w12_20,w12_21,w12_22,w12_23,w12_24,w12_25,w12_26,w12_27,w12_28,w12_29,w12_30,w12_31,w12_32,
		w12_33,w12_34,w12_35,w12_36,w12_37,w12_38,w12_39,w12_40,w12_41,w12_42,w12_43,w12_44,w12_45,w12_46,w12_47,w12_48,
		w12_49,w12_50,w12_51,w12_52,w12_53,w12_54,w12_55,w12_56,w12_57,w12_58,w12_59,w12_60,w12_61,w12_62,w12_63,w12_64,
		w12_65,w12_66,w12_67,w12_68,w12_69,w12_70,w12_71,w12_72,w12_73,w12_74,w12_75,w12_76,w12_77,w12_78,w12_79,w12_80,
		w12_81,w12_82,w12_83,w12_84,w12_85,w12_86,w12_87,w12_88,w12_89,w12_90,w12_91,w12_92,w12_93,w12_94,w12_95,w12_96,
		w12_97,w12_98,w12_99,w12_100,w12_101,w12_102,w12_103,w12_104,w12_105,w12_106,w12_107,w12_108,w12_109,w12_110,w12_111,w12_112,
		w12_113,w12_114,w12_115,w12_116,w12_117,w12_118,w12_119,w12_120,w12_121,w12_122,w12_123,w12_124,w12_125,w12_126,
	w13_0,w13_1,w13_2,w13_3,w13_4,w13_5,w13_6,w13_7,w13_8,w13_9,w13_10,w13_11,w13_12,w13_13,w13_14,w13_15,w13_16,
		w13_17,w13_18,w13_19,w13_20,w13_21,w13_22,w13_23,w13_24,w13_25,w13_26,w13_27,w13_28,w13_29,w13_30,w13_31,w13_32,
		w13_33,w13_34,w13_35,w13_36,w13_37,w13_38,w13_39,w13_40,w13_41,w13_42,w13_43,w13_44,w13_45,w13_46,w13_47,w13_48,
		w13_49,w13_50,w13_51,w13_52,w13_53,w13_54,w13_55,w13_56,w13_57,w13_58,w13_59,w13_60,w13_61,w13_62,w13_63,w13_64,
		w13_65,w13_66,w13_67,w13_68,w13_69,w13_70,w13_71,w13_72,w13_73,w13_74,w13_75,w13_76,w13_77,w13_78,w13_79,w13_80,
		w13_81,w13_82,w13_83,w13_84,w13_85,w13_86,w13_87,w13_88,w13_89,w13_90,w13_91,w13_92,w13_93,w13_94,w13_95,w13_96,
		w13_97,w13_98,w13_99,w13_100,w13_101,w13_102,w13_103,w13_104,w13_105,w13_106,w13_107,w13_108,w13_109,w13_110,w13_111,w13_112,
		w13_113,w13_114,w13_115,w13_116,w13_117,w13_118,w13_119,w13_120,w13_121,w13_122,w13_123,w13_124,w13_125,w13_126,
	w14_0,w14_1,w14_2,w14_3,w14_4,w14_5,w14_6,w14_7,w14_8,w14_9,w14_10,w14_11,w14_12,w14_13,w14_14,w14_15,w14_16,
		w14_17,w14_18,w14_19,w14_20,w14_21,w14_22,w14_23,w14_24,w14_25,w14_26,w14_27,w14_28,w14_29,w14_30,w14_31,w14_32,
		w14_33,w14_34,w14_35,w14_36,w14_37,w14_38,w14_39,w14_40,w14_41,w14_42,w14_43,w14_44,w14_45,w14_46,w14_47,w14_48,
		w14_49,w14_50,w14_51,w14_52,w14_53,w14_54,w14_55,w14_56,w14_57,w14_58,w14_59,w14_60,w14_61,w14_62,w14_63,w14_64,
		w14_65,w14_66,w14_67,w14_68,w14_69,w14_70,w14_71,w14_72,w14_73,w14_74,w14_75,w14_76,w14_77,w14_78,w14_79,w14_80,
		w14_81,w14_82,w14_83,w14_84,w14_85,w14_86,w14_87,w14_88,w14_89,w14_90,w14_91,w14_92,w14_93,w14_94,w14_95,w14_96,
		w14_97,w14_98,w14_99,w14_100,w14_101,w14_102,w14_103,w14_104,w14_105,w14_106,w14_107,w14_108,w14_109,w14_110,w14_111,w14_112,
		w14_113,w14_114,w14_115,w14_116,w14_117,w14_118,w14_119,w14_120,w14_121,w14_122,w14_123,w14_124,w14_125,w14_126,
	w15_0,w15_1,w15_2,w15_3,w15_4,w15_5,w15_6,w15_7,w15_8,w15_9,w15_10,w15_11,w15_12,w15_13,w15_14,w15_15,w15_16,
		w15_17,w15_18,w15_19,w15_20,w15_21,w15_22,w15_23,w15_24,w15_25,w15_26,w15_27,w15_28,w15_29,w15_30,w15_31,w15_32,
		w15_33,w15_34,w15_35,w15_36,w15_37,w15_38,w15_39,w15_40,w15_41,w15_42,w15_43,w15_44,w15_45,w15_46,w15_47,w15_48,
		w15_49,w15_50,w15_51,w15_52,w15_53,w15_54,w15_55,w15_56,w15_57,w15_58,w15_59,w15_60,w15_61,w15_62,w15_63,w15_64,
		w15_65,w15_66,w15_67,w15_68,w15_69,w15_70,w15_71,w15_72,w15_73,w15_74,w15_75,w15_76,w15_77,w15_78,w15_79,w15_80,
		w15_81,w15_82,w15_83,w15_84,w15_85,w15_86,w15_87,w15_88,w15_89,w15_90,w15_91,w15_92,w15_93,w15_94,w15_95,w15_96,
		w15_97,w15_98,w15_99,w15_100,w15_101,w15_102,w15_103,w15_104,w15_105,w15_106,w15_107,w15_108,w15_109,w15_110,w15_111,w15_112,
		w15_113,w15_114,w15_115,w15_116,w15_117,w15_118,w15_119,w15_120,w15_121,w15_122,w15_123,w15_124,w15_125,w15_126,
	w16_0,w16_1,w16_2,w16_3,w16_4,w16_5,w16_6,w16_7,w16_8,w16_9,w16_10,w16_11,w16_12,w16_13,w16_14,w16_15,w16_16,
		w16_17,w16_18,w16_19,w16_20,w16_21,w16_22,w16_23,w16_24,w16_25,w16_26,w16_27,w16_28,w16_29,w16_30,w16_31,w16_32,
		w16_33,w16_34,w16_35,w16_36,w16_37,w16_38,w16_39,w16_40,w16_41,w16_42,w16_43,w16_44,w16_45,w16_46,w16_47,w16_48,
		w16_49,w16_50,w16_51,w16_52,w16_53,w16_54,w16_55,w16_56,w16_57,w16_58,w16_59,w16_60,w16_61,w16_62,w16_63,w16_64,
		w16_65,w16_66,w16_67,w16_68,w16_69,w16_70,w16_71,w16_72,w16_73,w16_74,w16_75,w16_76,w16_77,w16_78,w16_79,w16_80,
		w16_81,w16_82,w16_83,w16_84,w16_85,w16_86,w16_87,w16_88,w16_89,w16_90,w16_91,w16_92,w16_93,w16_94,w16_95,w16_96,
		w16_97,w16_98,w16_99,w16_100,w16_101,w16_102,w16_103,w16_104,w16_105,w16_106,w16_107,w16_108,w16_109,w16_110,w16_111,w16_112,
		w16_113,w16_114,w16_115,w16_116,w16_117,w16_118,w16_119,w16_120,w16_121,w16_122,w16_123,w16_124,w16_125,w16_126,
	w17_0,w17_1,w17_2,w17_3,w17_4,w17_5,w17_6,w17_7,w17_8,w17_9,w17_10,w17_11,w17_12,w17_13,w17_14,w17_15,w17_16,
		w17_17,w17_18,w17_19,w17_20,w17_21,w17_22,w17_23,w17_24,w17_25,w17_26,w17_27,w17_28,w17_29,w17_30,w17_31,w17_32,
		w17_33,w17_34,w17_35,w17_36,w17_37,w17_38,w17_39,w17_40,w17_41,w17_42,w17_43,w17_44,w17_45,w17_46,w17_47,w17_48,
		w17_49,w17_50,w17_51,w17_52,w17_53,w17_54,w17_55,w17_56,w17_57,w17_58,w17_59,w17_60,w17_61,w17_62,w17_63,w17_64,
		w17_65,w17_66,w17_67,w17_68,w17_69,w17_70,w17_71,w17_72,w17_73,w17_74,w17_75,w17_76,w17_77,w17_78,w17_79,w17_80,
		w17_81,w17_82,w17_83,w17_84,w17_85,w17_86,w17_87,w17_88,w17_89,w17_90,w17_91,w17_92,w17_93,w17_94,w17_95,w17_96,
		w17_97,w17_98,w17_99,w17_100,w17_101,w17_102,w17_103,w17_104,w17_105,w17_106,w17_107,w17_108,w17_109,w17_110,w17_111,w17_112,
		w17_113,w17_114,w17_115,w17_116,w17_117,w17_118,w17_119,w17_120,w17_121,w17_122,w17_123,w17_124,w17_125,w17_126,
	w18_0,w18_1,w18_2,w18_3,w18_4,w18_5,w18_6,w18_7,w18_8,w18_9,w18_10,w18_11,w18_12,w18_13,w18_14,w18_15,w18_16,
		w18_17,w18_18,w18_19,w18_20,w18_21,w18_22,w18_23,w18_24,w18_25,w18_26,w18_27,w18_28,w18_29,w18_30,w18_31,w18_32,
		w18_33,w18_34,w18_35,w18_36,w18_37,w18_38,w18_39,w18_40,w18_41,w18_42,w18_43,w18_44,w18_45,w18_46,w18_47,w18_48,
		w18_49,w18_50,w18_51,w18_52,w18_53,w18_54,w18_55,w18_56,w18_57,w18_58,w18_59,w18_60,w18_61,w18_62,w18_63,w18_64,
		w18_65,w18_66,w18_67,w18_68,w18_69,w18_70,w18_71,w18_72,w18_73,w18_74,w18_75,w18_76,w18_77,w18_78,w18_79,w18_80,
		w18_81,w18_82,w18_83,w18_84,w18_85,w18_86,w18_87,w18_88,w18_89,w18_90,w18_91,w18_92,w18_93,w18_94,w18_95,w18_96,
		w18_97,w18_98,w18_99,w18_100,w18_101,w18_102,w18_103,w18_104,w18_105,w18_106,w18_107,w18_108,w18_109,w18_110,w18_111,w18_112,
		w18_113,w18_114,w18_115,w18_116,w18_117,w18_118,w18_119,w18_120,w18_121,w18_122,w18_123,w18_124,w18_125,w18_126,
	w19_0,w19_1,w19_2,w19_3,w19_4,w19_5,w19_6,w19_7,w19_8,w19_9,w19_10,w19_11,w19_12,w19_13,w19_14,w19_15,w19_16,
		w19_17,w19_18,w19_19,w19_20,w19_21,w19_22,w19_23,w19_24,w19_25,w19_26,w19_27,w19_28,w19_29,w19_30,w19_31,w19_32,
		w19_33,w19_34,w19_35,w19_36,w19_37,w19_38,w19_39,w19_40,w19_41,w19_42,w19_43,w19_44,w19_45,w19_46,w19_47,w19_48,
		w19_49,w19_50,w19_51,w19_52,w19_53,w19_54,w19_55,w19_56,w19_57,w19_58,w19_59,w19_60,w19_61,w19_62,w19_63,w19_64,
		w19_65,w19_66,w19_67,w19_68,w19_69,w19_70,w19_71,w19_72,w19_73,w19_74,w19_75,w19_76,w19_77,w19_78,w19_79,w19_80,
		w19_81,w19_82,w19_83,w19_84,w19_85,w19_86,w19_87,w19_88,w19_89,w19_90,w19_91,w19_92,w19_93,w19_94,w19_95,w19_96,
		w19_97,w19_98,w19_99,w19_100,w19_101,w19_102,w19_103,w19_104,w19_105,w19_106,w19_107,w19_108,w19_109,w19_110,w19_111,w19_112,
		w19_113,w19_114,w19_115,w19_116,w19_117,w19_118,w19_119,w19_120,w19_121,w19_122,w19_123,w19_124,w19_125,w19_126,
	w20_0,w20_1,w20_2,w20_3,w20_4,w20_5,w20_6,w20_7,w20_8,w20_9,w20_10,w20_11,w20_12,w20_13,w20_14,w20_15,w20_16,
		w20_17,w20_18,w20_19,w20_20,w20_21,w20_22,w20_23,w20_24,w20_25,w20_26,w20_27,w20_28,w20_29,w20_30,w20_31,w20_32,
		w20_33,w20_34,w20_35,w20_36,w20_37,w20_38,w20_39,w20_40,w20_41,w20_42,w20_43,w20_44,w20_45,w20_46,w20_47,w20_48,
		w20_49,w20_50,w20_51,w20_52,w20_53,w20_54,w20_55,w20_56,w20_57,w20_58,w20_59,w20_60,w20_61,w20_62,w20_63,w20_64,
		w20_65,w20_66,w20_67,w20_68,w20_69,w20_70,w20_71,w20_72,w20_73,w20_74,w20_75,w20_76,w20_77,w20_78,w20_79,w20_80,
		w20_81,w20_82,w20_83,w20_84,w20_85,w20_86,w20_87,w20_88,w20_89,w20_90,w20_91,w20_92,w20_93,w20_94,w20_95,w20_96,
		w20_97,w20_98,w20_99,w20_100,w20_101,w20_102,w20_103,w20_104,w20_105,w20_106,w20_107,w20_108,w20_109,w20_110,w20_111,w20_112,
		w20_113,w20_114,w20_115,w20_116,w20_117,w20_118,w20_119,w20_120,w20_121,w20_122,w20_123,w20_124,w20_125,w20_126,
	w21_0,w21_1,w21_2,w21_3,w21_4,w21_5,w21_6,w21_7,w21_8,w21_9,w21_10,w21_11,w21_12,w21_13,w21_14,w21_15,w21_16,
		w21_17,w21_18,w21_19,w21_20,w21_21,w21_22,w21_23,w21_24,w21_25,w21_26,w21_27,w21_28,w21_29,w21_30,w21_31,w21_32,
		w21_33,w21_34,w21_35,w21_36,w21_37,w21_38,w21_39,w21_40,w21_41,w21_42,w21_43,w21_44,w21_45,w21_46,w21_47,w21_48,
		w21_49,w21_50,w21_51,w21_52,w21_53,w21_54,w21_55,w21_56,w21_57,w21_58,w21_59,w21_60,w21_61,w21_62,w21_63,w21_64,
		w21_65,w21_66,w21_67,w21_68,w21_69,w21_70,w21_71,w21_72,w21_73,w21_74,w21_75,w21_76,w21_77,w21_78,w21_79,w21_80,
		w21_81,w21_82,w21_83,w21_84,w21_85,w21_86,w21_87,w21_88,w21_89,w21_90,w21_91,w21_92,w21_93,w21_94,w21_95,w21_96,
		w21_97,w21_98,w21_99,w21_100,w21_101,w21_102,w21_103,w21_104,w21_105,w21_106,w21_107,w21_108,w21_109,w21_110,w21_111,w21_112,
		w21_113,w21_114,w21_115,w21_116,w21_117,w21_118,w21_119,w21_120,w21_121,w21_122,w21_123,w21_124,w21_125,w21_126,
	w22_0,w22_1,w22_2,w22_3,w22_4,w22_5,w22_6,w22_7,w22_8,w22_9,w22_10,w22_11,w22_12,w22_13,w22_14,w22_15,w22_16,
		w22_17,w22_18,w22_19,w22_20,w22_21,w22_22,w22_23,w22_24,w22_25,w22_26,w22_27,w22_28,w22_29,w22_30,w22_31,w22_32,
		w22_33,w22_34,w22_35,w22_36,w22_37,w22_38,w22_39,w22_40,w22_41,w22_42,w22_43,w22_44,w22_45,w22_46,w22_47,w22_48,
		w22_49,w22_50,w22_51,w22_52,w22_53,w22_54,w22_55,w22_56,w22_57,w22_58,w22_59,w22_60,w22_61,w22_62,w22_63,w22_64,
		w22_65,w22_66,w22_67,w22_68,w22_69,w22_70,w22_71,w22_72,w22_73,w22_74,w22_75,w22_76,w22_77,w22_78,w22_79,w22_80,
		w22_81,w22_82,w22_83,w22_84,w22_85,w22_86,w22_87,w22_88,w22_89,w22_90,w22_91,w22_92,w22_93,w22_94,w22_95,w22_96,
		w22_97,w22_98,w22_99,w22_100,w22_101,w22_102,w22_103,w22_104,w22_105,w22_106,w22_107,w22_108,w22_109,w22_110,w22_111,w22_112,
		w22_113,w22_114,w22_115,w22_116,w22_117,w22_118,w22_119,w22_120,w22_121,w22_122,w22_123,w22_124,w22_125,w22_126,
	w23_0,w23_1,w23_2,w23_3,w23_4,w23_5,w23_6,w23_7,w23_8,w23_9,w23_10,w23_11,w23_12,w23_13,w23_14,w23_15,w23_16,
		w23_17,w23_18,w23_19,w23_20,w23_21,w23_22,w23_23,w23_24,w23_25,w23_26,w23_27,w23_28,w23_29,w23_30,w23_31,w23_32,
		w23_33,w23_34,w23_35,w23_36,w23_37,w23_38,w23_39,w23_40,w23_41,w23_42,w23_43,w23_44,w23_45,w23_46,w23_47,w23_48,
		w23_49,w23_50,w23_51,w23_52,w23_53,w23_54,w23_55,w23_56,w23_57,w23_58,w23_59,w23_60,w23_61,w23_62,w23_63,w23_64,
		w23_65,w23_66,w23_67,w23_68,w23_69,w23_70,w23_71,w23_72,w23_73,w23_74,w23_75,w23_76,w23_77,w23_78,w23_79,w23_80,
		w23_81,w23_82,w23_83,w23_84,w23_85,w23_86,w23_87,w23_88,w23_89,w23_90,w23_91,w23_92,w23_93,w23_94,w23_95,w23_96,
		w23_97,w23_98,w23_99,w23_100,w23_101,w23_102,w23_103,w23_104,w23_105,w23_106,w23_107,w23_108,w23_109,w23_110,w23_111,w23_112,
		w23_113,w23_114,w23_115,w23_116,w23_117,w23_118,w23_119,w23_120,w23_121,w23_122,w23_123,w23_124,w23_125,w23_126,
	w24_0,w24_1,w24_2,w24_3,w24_4,w24_5,w24_6,w24_7,w24_8,w24_9,w24_10,w24_11,w24_12,w24_13,w24_14,w24_15,w24_16,
		w24_17,w24_18,w24_19,w24_20,w24_21,w24_22,w24_23,w24_24,w24_25,w24_26,w24_27,w24_28,w24_29,w24_30,w24_31,w24_32,
		w24_33,w24_34,w24_35,w24_36,w24_37,w24_38,w24_39,w24_40,w24_41,w24_42,w24_43,w24_44,w24_45,w24_46,w24_47,w24_48,
		w24_49,w24_50,w24_51,w24_52,w24_53,w24_54,w24_55,w24_56,w24_57,w24_58,w24_59,w24_60,w24_61,w24_62,w24_63,w24_64,
		w24_65,w24_66,w24_67,w24_68,w24_69,w24_70,w24_71,w24_72,w24_73,w24_74,w24_75,w24_76,w24_77,w24_78,w24_79,w24_80,
		w24_81,w24_82,w24_83,w24_84,w24_85,w24_86,w24_87,w24_88,w24_89,w24_90,w24_91,w24_92,w24_93,w24_94,w24_95,w24_96,
		w24_97,w24_98,w24_99,w24_100,w24_101,w24_102,w24_103,w24_104,w24_105,w24_106,w24_107,w24_108,w24_109,w24_110,w24_111,w24_112,
		w24_113,w24_114,w24_115,w24_116,w24_117,w24_118,w24_119,w24_120,w24_121,w24_122,w24_123,w24_124,w24_125,w24_126,
	w25_0,w25_1,w25_2,w25_3,w25_4,w25_5,w25_6,w25_7,w25_8,w25_9,w25_10,w25_11,w25_12,w25_13,w25_14,w25_15,w25_16,
		w25_17,w25_18,w25_19,w25_20,w25_21,w25_22,w25_23,w25_24,w25_25,w25_26,w25_27,w25_28,w25_29,w25_30,w25_31,w25_32,
		w25_33,w25_34,w25_35,w25_36,w25_37,w25_38,w25_39,w25_40,w25_41,w25_42,w25_43,w25_44,w25_45,w25_46,w25_47,w25_48,
		w25_49,w25_50,w25_51,w25_52,w25_53,w25_54,w25_55,w25_56,w25_57,w25_58,w25_59,w25_60,w25_61,w25_62,w25_63,w25_64,
		w25_65,w25_66,w25_67,w25_68,w25_69,w25_70,w25_71,w25_72,w25_73,w25_74,w25_75,w25_76,w25_77,w25_78,w25_79,w25_80,
		w25_81,w25_82,w25_83,w25_84,w25_85,w25_86,w25_87,w25_88,w25_89,w25_90,w25_91,w25_92,w25_93,w25_94,w25_95,w25_96,
		w25_97,w25_98,w25_99,w25_100,w25_101,w25_102,w25_103,w25_104,w25_105,w25_106,w25_107,w25_108,w25_109,w25_110,w25_111,w25_112,
		w25_113,w25_114,w25_115,w25_116,w25_117,w25_118,w25_119,w25_120,w25_121,w25_122,w25_123,w25_124,w25_125,w25_126,
	w26_0,w26_1,w26_2,w26_3,w26_4,w26_5,w26_6,w26_7,w26_8,w26_9,w26_10,w26_11,w26_12,w26_13,w26_14,w26_15,w26_16,
		w26_17,w26_18,w26_19,w26_20,w26_21,w26_22,w26_23,w26_24,w26_25,w26_26,w26_27,w26_28,w26_29,w26_30,w26_31,w26_32,
		w26_33,w26_34,w26_35,w26_36,w26_37,w26_38,w26_39,w26_40,w26_41,w26_42,w26_43,w26_44,w26_45,w26_46,w26_47,w26_48,
		w26_49,w26_50,w26_51,w26_52,w26_53,w26_54,w26_55,w26_56,w26_57,w26_58,w26_59,w26_60,w26_61,w26_62,w26_63,w26_64,
		w26_65,w26_66,w26_67,w26_68,w26_69,w26_70,w26_71,w26_72,w26_73,w26_74,w26_75,w26_76,w26_77,w26_78,w26_79,w26_80,
		w26_81,w26_82,w26_83,w26_84,w26_85,w26_86,w26_87,w26_88,w26_89,w26_90,w26_91,w26_92,w26_93,w26_94,w26_95,w26_96,
		w26_97,w26_98,w26_99,w26_100,w26_101,w26_102,w26_103,w26_104,w26_105,w26_106,w26_107,w26_108,w26_109,w26_110,w26_111,w26_112,
		w26_113,w26_114,w26_115,w26_116,w26_117,w26_118,w26_119,w26_120,w26_121,w26_122,w26_123,w26_124,w26_125,w26_126,
	w27_0,w27_1,w27_2,w27_3,w27_4,w27_5,w27_6,w27_7,w27_8,w27_9,w27_10,w27_11,w27_12,w27_13,w27_14,w27_15,w27_16,
		w27_17,w27_18,w27_19,w27_20,w27_21,w27_22,w27_23,w27_24,w27_25,w27_26,w27_27,w27_28,w27_29,w27_30,w27_31,w27_32,
		w27_33,w27_34,w27_35,w27_36,w27_37,w27_38,w27_39,w27_40,w27_41,w27_42,w27_43,w27_44,w27_45,w27_46,w27_47,w27_48,
		w27_49,w27_50,w27_51,w27_52,w27_53,w27_54,w27_55,w27_56,w27_57,w27_58,w27_59,w27_60,w27_61,w27_62,w27_63,w27_64,
		w27_65,w27_66,w27_67,w27_68,w27_69,w27_70,w27_71,w27_72,w27_73,w27_74,w27_75,w27_76,w27_77,w27_78,w27_79,w27_80,
		w27_81,w27_82,w27_83,w27_84,w27_85,w27_86,w27_87,w27_88,w27_89,w27_90,w27_91,w27_92,w27_93,w27_94,w27_95,w27_96,
		w27_97,w27_98,w27_99,w27_100,w27_101,w27_102,w27_103,w27_104,w27_105,w27_106,w27_107,w27_108,w27_109,w27_110,w27_111,w27_112,
		w27_113,w27_114,w27_115,w27_116,w27_117,w27_118,w27_119,w27_120,w27_121,w27_122,w27_123,w27_124,w27_125,w27_126,
	w28_0,w28_1,w28_2,w28_3,w28_4,w28_5,w28_6,w28_7,w28_8,w28_9,w28_10,w28_11,w28_12,w28_13,w28_14,w28_15,w28_16,
		w28_17,w28_18,w28_19,w28_20,w28_21,w28_22,w28_23,w28_24,w28_25,w28_26,w28_27,w28_28,w28_29,w28_30,w28_31,w28_32,
		w28_33,w28_34,w28_35,w28_36,w28_37,w28_38,w28_39,w28_40,w28_41,w28_42,w28_43,w28_44,w28_45,w28_46,w28_47,w28_48,
		w28_49,w28_50,w28_51,w28_52,w28_53,w28_54,w28_55,w28_56,w28_57,w28_58,w28_59,w28_60,w28_61,w28_62,w28_63,w28_64,
		w28_65,w28_66,w28_67,w28_68,w28_69,w28_70,w28_71,w28_72,w28_73,w28_74,w28_75,w28_76,w28_77,w28_78,w28_79,w28_80,
		w28_81,w28_82,w28_83,w28_84,w28_85,w28_86,w28_87,w28_88,w28_89,w28_90,w28_91,w28_92,w28_93,w28_94,w28_95,w28_96,
		w28_97,w28_98,w28_99,w28_100,w28_101,w28_102,w28_103,w28_104,w28_105,w28_106,w28_107,w28_108,w28_109,w28_110,w28_111,w28_112,
		w28_113,w28_114,w28_115,w28_116,w28_117,w28_118,w28_119,w28_120,w28_121,w28_122,w28_123,w28_124,w28_125,w28_126,
	w29_0,w29_1,w29_2,w29_3,w29_4,w29_5,w29_6,w29_7,w29_8,w29_9,w29_10,w29_11,w29_12,w29_13,w29_14,w29_15,w29_16,
		w29_17,w29_18,w29_19,w29_20,w29_21,w29_22,w29_23,w29_24,w29_25,w29_26,w29_27,w29_28,w29_29,w29_30,w29_31,w29_32,
		w29_33,w29_34,w29_35,w29_36,w29_37,w29_38,w29_39,w29_40,w29_41,w29_42,w29_43,w29_44,w29_45,w29_46,w29_47,w29_48,
		w29_49,w29_50,w29_51,w29_52,w29_53,w29_54,w29_55,w29_56,w29_57,w29_58,w29_59,w29_60,w29_61,w29_62,w29_63,w29_64,
		w29_65,w29_66,w29_67,w29_68,w29_69,w29_70,w29_71,w29_72,w29_73,w29_74,w29_75,w29_76,w29_77,w29_78,w29_79,w29_80,
		w29_81,w29_82,w29_83,w29_84,w29_85,w29_86,w29_87,w29_88,w29_89,w29_90,w29_91,w29_92,w29_93,w29_94,w29_95,w29_96,
		w29_97,w29_98,w29_99,w29_100,w29_101,w29_102,w29_103,w29_104,w29_105,w29_106,w29_107,w29_108,w29_109,w29_110,w29_111,w29_112,
		w29_113,w29_114,w29_115,w29_116,w29_117,w29_118,w29_119,w29_120,w29_121,w29_122,w29_123,w29_124,w29_125,w29_126,
	w30_0,w30_1,w30_2,w30_3,w30_4,w30_5,w30_6,w30_7,w30_8,w30_9,w30_10,w30_11,w30_12,w30_13,w30_14,w30_15,w30_16,
		w30_17,w30_18,w30_19,w30_20,w30_21,w30_22,w30_23,w30_24,w30_25,w30_26,w30_27,w30_28,w30_29,w30_30,w30_31,w30_32,
		w30_33,w30_34,w30_35,w30_36,w30_37,w30_38,w30_39,w30_40,w30_41,w30_42,w30_43,w30_44,w30_45,w30_46,w30_47,w30_48,
		w30_49,w30_50,w30_51,w30_52,w30_53,w30_54,w30_55,w30_56,w30_57,w30_58,w30_59,w30_60,w30_61,w30_62,w30_63,w30_64,
		w30_65,w30_66,w30_67,w30_68,w30_69,w30_70,w30_71,w30_72,w30_73,w30_74,w30_75,w30_76,w30_77,w30_78,w30_79,w30_80,
		w30_81,w30_82,w30_83,w30_84,w30_85,w30_86,w30_87,w30_88,w30_89,w30_90,w30_91,w30_92,w30_93,w30_94,w30_95,w30_96,
		w30_97,w30_98,w30_99,w30_100,w30_101,w30_102,w30_103,w30_104,w30_105,w30_106,w30_107,w30_108,w30_109,w30_110,w30_111,w30_112,
		w30_113,w30_114,w30_115,w30_116,w30_117,w30_118,w30_119,w30_120,w30_121,w30_122,w30_123,w30_124,w30_125,w30_126,
	w31_0,w31_1,w31_2,w31_3,w31_4,w31_5,w31_6,w31_7,w31_8,w31_9,w31_10,w31_11,w31_12,w31_13,w31_14,w31_15,w31_16,
		w31_17,w31_18,w31_19,w31_20,w31_21,w31_22,w31_23,w31_24,w31_25,w31_26,w31_27,w31_28,w31_29,w31_30,w31_31,w31_32,
		w31_33,w31_34,w31_35,w31_36,w31_37,w31_38,w31_39,w31_40,w31_41,w31_42,w31_43,w31_44,w31_45,w31_46,w31_47,w31_48,
		w31_49,w31_50,w31_51,w31_52,w31_53,w31_54,w31_55,w31_56,w31_57,w31_58,w31_59,w31_60,w31_61,w31_62,w31_63,w31_64,
		w31_65,w31_66,w31_67,w31_68,w31_69,w31_70,w31_71,w31_72,w31_73,w31_74,w31_75,w31_76,w31_77,w31_78,w31_79,w31_80,
		w31_81,w31_82,w31_83,w31_84,w31_85,w31_86,w31_87,w31_88,w31_89,w31_90,w31_91,w31_92,w31_93,w31_94,w31_95,w31_96,
		w31_97,w31_98,w31_99,w31_100,w31_101,w31_102,w31_103,w31_104,w31_105,w31_106,w31_107,w31_108,w31_109,w31_110,w31_111,w31_112,
		w31_113,w31_114,w31_115,w31_116,w31_117,w31_118,w31_119,w31_120,w31_121,w31_122,w31_123,w31_124,w31_125,w31_126,
	w32_0,w32_1,w32_2,w32_3,w32_4,w32_5,w32_6,w32_7,w32_8,w32_9,w32_10,w32_11,w32_12,w32_13,w32_14,w32_15,w32_16,
		w32_17,w32_18,w32_19,w32_20,w32_21,w32_22,w32_23,w32_24,w32_25,w32_26,w32_27,w32_28,w32_29,w32_30,w32_31,w32_32,
		w32_33,w32_34,w32_35,w32_36,w32_37,w32_38,w32_39,w32_40,w32_41,w32_42,w32_43,w32_44,w32_45,w32_46,w32_47,w32_48,
		w32_49,w32_50,w32_51,w32_52,w32_53,w32_54,w32_55,w32_56,w32_57,w32_58,w32_59,w32_60,w32_61,w32_62,w32_63,w32_64,
		w32_65,w32_66,w32_67,w32_68,w32_69,w32_70,w32_71,w32_72,w32_73,w32_74,w32_75,w32_76,w32_77,w32_78,w32_79,w32_80,
		w32_81,w32_82,w32_83,w32_84,w32_85,w32_86,w32_87,w32_88,w32_89,w32_90,w32_91,w32_92,w32_93,w32_94,w32_95,w32_96,
		w32_97,w32_98,w32_99,w32_100,w32_101,w32_102,w32_103,w32_104,w32_105,w32_106,w32_107,w32_108,w32_109,w32_110,w32_111,w32_112,
		w32_113,w32_114,w32_115,w32_116,w32_117,w32_118,w32_119,w32_120,w32_121,w32_122,w32_123,w32_124,w32_125,w32_126,
	w33_0,w33_1,w33_2,w33_3,w33_4,w33_5,w33_6,w33_7,w33_8,w33_9,w33_10,w33_11,w33_12,w33_13,w33_14,w33_15,w33_16,
		w33_17,w33_18,w33_19,w33_20,w33_21,w33_22,w33_23,w33_24,w33_25,w33_26,w33_27,w33_28,w33_29,w33_30,w33_31,w33_32,
		w33_33,w33_34,w33_35,w33_36,w33_37,w33_38,w33_39,w33_40,w33_41,w33_42,w33_43,w33_44,w33_45,w33_46,w33_47,w33_48,
		w33_49,w33_50,w33_51,w33_52,w33_53,w33_54,w33_55,w33_56,w33_57,w33_58,w33_59,w33_60,w33_61,w33_62,w33_63,w33_64,
		w33_65,w33_66,w33_67,w33_68,w33_69,w33_70,w33_71,w33_72,w33_73,w33_74,w33_75,w33_76,w33_77,w33_78,w33_79,w33_80,
		w33_81,w33_82,w33_83,w33_84,w33_85,w33_86,w33_87,w33_88,w33_89,w33_90,w33_91,w33_92,w33_93,w33_94,w33_95,w33_96,
		w33_97,w33_98,w33_99,w33_100,w33_101,w33_102,w33_103,w33_104,w33_105,w33_106,w33_107,w33_108,w33_109,w33_110,w33_111,w33_112,
		w33_113,w33_114,w33_115,w33_116,w33_117,w33_118,w33_119,w33_120,w33_121,w33_122,w33_123,w33_124,w33_125,w33_126,
	w34_0,w34_1,w34_2,w34_3,w34_4,w34_5,w34_6,w34_7,w34_8,w34_9,w34_10,w34_11,w34_12,w34_13,w34_14,w34_15,w34_16,
		w34_17,w34_18,w34_19,w34_20,w34_21,w34_22,w34_23,w34_24,w34_25,w34_26,w34_27,w34_28,w34_29,w34_30,w34_31,w34_32,
		w34_33,w34_34,w34_35,w34_36,w34_37,w34_38,w34_39,w34_40,w34_41,w34_42,w34_43,w34_44,w34_45,w34_46,w34_47,w34_48,
		w34_49,w34_50,w34_51,w34_52,w34_53,w34_54,w34_55,w34_56,w34_57,w34_58,w34_59,w34_60,w34_61,w34_62,w34_63,w34_64,
		w34_65,w34_66,w34_67,w34_68,w34_69,w34_70,w34_71,w34_72,w34_73,w34_74,w34_75,w34_76,w34_77,w34_78,w34_79,w34_80,
		w34_81,w34_82,w34_83,w34_84,w34_85,w34_86,w34_87,w34_88,w34_89,w34_90,w34_91,w34_92,w34_93,w34_94,w34_95,w34_96,
		w34_97,w34_98,w34_99,w34_100,w34_101,w34_102,w34_103,w34_104,w34_105,w34_106,w34_107,w34_108,w34_109,w34_110,w34_111,w34_112,
		w34_113,w34_114,w34_115,w34_116,w34_117,w34_118,w34_119,w34_120,w34_121,w34_122,w34_123,w34_124,w34_125,w34_126,
	w35_0,w35_1,w35_2,w35_3,w35_4,w35_5,w35_6,w35_7,w35_8,w35_9,w35_10,w35_11,w35_12,w35_13,w35_14,w35_15,w35_16,
		w35_17,w35_18,w35_19,w35_20,w35_21,w35_22,w35_23,w35_24,w35_25,w35_26,w35_27,w35_28,w35_29,w35_30,w35_31,w35_32,
		w35_33,w35_34,w35_35,w35_36,w35_37,w35_38,w35_39,w35_40,w35_41,w35_42,w35_43,w35_44,w35_45,w35_46,w35_47,w35_48,
		w35_49,w35_50,w35_51,w35_52,w35_53,w35_54,w35_55,w35_56,w35_57,w35_58,w35_59,w35_60,w35_61,w35_62,w35_63,w35_64,
		w35_65,w35_66,w35_67,w35_68,w35_69,w35_70,w35_71,w35_72,w35_73,w35_74,w35_75,w35_76,w35_77,w35_78,w35_79,w35_80,
		w35_81,w35_82,w35_83,w35_84,w35_85,w35_86,w35_87,w35_88,w35_89,w35_90,w35_91,w35_92,w35_93,w35_94,w35_95,w35_96,
		w35_97,w35_98,w35_99,w35_100,w35_101,w35_102,w35_103,w35_104,w35_105,w35_106,w35_107,w35_108,w35_109,w35_110,w35_111,w35_112,
		w35_113,w35_114,w35_115,w35_116,w35_117,w35_118,w35_119,w35_120,w35_121,w35_122,w35_123,w35_124,w35_125,w35_126,
	w36_0,w36_1,w36_2,w36_3,w36_4,w36_5,w36_6,w36_7,w36_8,w36_9,w36_10,w36_11,w36_12,w36_13,w36_14,w36_15,w36_16,
		w36_17,w36_18,w36_19,w36_20,w36_21,w36_22,w36_23,w36_24,w36_25,w36_26,w36_27,w36_28,w36_29,w36_30,w36_31,w36_32,
		w36_33,w36_34,w36_35,w36_36,w36_37,w36_38,w36_39,w36_40,w36_41,w36_42,w36_43,w36_44,w36_45,w36_46,w36_47,w36_48,
		w36_49,w36_50,w36_51,w36_52,w36_53,w36_54,w36_55,w36_56,w36_57,w36_58,w36_59,w36_60,w36_61,w36_62,w36_63,w36_64,
		w36_65,w36_66,w36_67,w36_68,w36_69,w36_70,w36_71,w36_72,w36_73,w36_74,w36_75,w36_76,w36_77,w36_78,w36_79,w36_80,
		w36_81,w36_82,w36_83,w36_84,w36_85,w36_86,w36_87,w36_88,w36_89,w36_90,w36_91,w36_92,w36_93,w36_94,w36_95,w36_96,
		w36_97,w36_98,w36_99,w36_100,w36_101,w36_102,w36_103,w36_104,w36_105,w36_106,w36_107,w36_108,w36_109,w36_110,w36_111,w36_112,
		w36_113,w36_114,w36_115,w36_116,w36_117,w36_118,w36_119,w36_120,w36_121,w36_122,w36_123,w36_124,w36_125,w36_126,
	w37_0,w37_1,w37_2,w37_3,w37_4,w37_5,w37_6,w37_7,w37_8,w37_9,w37_10,w37_11,w37_12,w37_13,w37_14,w37_15,w37_16,
		w37_17,w37_18,w37_19,w37_20,w37_21,w37_22,w37_23,w37_24,w37_25,w37_26,w37_27,w37_28,w37_29,w37_30,w37_31,w37_32,
		w37_33,w37_34,w37_35,w37_36,w37_37,w37_38,w37_39,w37_40,w37_41,w37_42,w37_43,w37_44,w37_45,w37_46,w37_47,w37_48,
		w37_49,w37_50,w37_51,w37_52,w37_53,w37_54,w37_55,w37_56,w37_57,w37_58,w37_59,w37_60,w37_61,w37_62,w37_63,w37_64,
		w37_65,w37_66,w37_67,w37_68,w37_69,w37_70,w37_71,w37_72,w37_73,w37_74,w37_75,w37_76,w37_77,w37_78,w37_79,w37_80,
		w37_81,w37_82,w37_83,w37_84,w37_85,w37_86,w37_87,w37_88,w37_89,w37_90,w37_91,w37_92,w37_93,w37_94,w37_95,w37_96,
		w37_97,w37_98,w37_99,w37_100,w37_101,w37_102,w37_103,w37_104,w37_105,w37_106,w37_107,w37_108,w37_109,w37_110,w37_111,w37_112,
		w37_113,w37_114,w37_115,w37_116,w37_117,w37_118,w37_119,w37_120,w37_121,w37_122,w37_123,w37_124,w37_125,w37_126,
	w38_0,w38_1,w38_2,w38_3,w38_4,w38_5,w38_6,w38_7,w38_8,w38_9,w38_10,w38_11,w38_12,w38_13,w38_14,w38_15,w38_16,
		w38_17,w38_18,w38_19,w38_20,w38_21,w38_22,w38_23,w38_24,w38_25,w38_26,w38_27,w38_28,w38_29,w38_30,w38_31,w38_32,
		w38_33,w38_34,w38_35,w38_36,w38_37,w38_38,w38_39,w38_40,w38_41,w38_42,w38_43,w38_44,w38_45,w38_46,w38_47,w38_48,
		w38_49,w38_50,w38_51,w38_52,w38_53,w38_54,w38_55,w38_56,w38_57,w38_58,w38_59,w38_60,w38_61,w38_62,w38_63,w38_64,
		w38_65,w38_66,w38_67,w38_68,w38_69,w38_70,w38_71,w38_72,w38_73,w38_74,w38_75,w38_76,w38_77,w38_78,w38_79,w38_80,
		w38_81,w38_82,w38_83,w38_84,w38_85,w38_86,w38_87,w38_88,w38_89,w38_90,w38_91,w38_92,w38_93,w38_94,w38_95,w38_96,
		w38_97,w38_98,w38_99,w38_100,w38_101,w38_102,w38_103,w38_104,w38_105,w38_106,w38_107,w38_108,w38_109,w38_110,w38_111,w38_112,
		w38_113,w38_114,w38_115,w38_116,w38_117,w38_118,w38_119,w38_120,w38_121,w38_122,w38_123,w38_124,w38_125,w38_126,
	w39_0,w39_1,w39_2,w39_3,w39_4,w39_5,w39_6,w39_7,w39_8,w39_9,w39_10,w39_11,w39_12,w39_13,w39_14,w39_15,w39_16,
		w39_17,w39_18,w39_19,w39_20,w39_21,w39_22,w39_23,w39_24,w39_25,w39_26,w39_27,w39_28,w39_29,w39_30,w39_31,w39_32,
		w39_33,w39_34,w39_35,w39_36,w39_37,w39_38,w39_39,w39_40,w39_41,w39_42,w39_43,w39_44,w39_45,w39_46,w39_47,w39_48,
		w39_49,w39_50,w39_51,w39_52,w39_53,w39_54,w39_55,w39_56,w39_57,w39_58,w39_59,w39_60,w39_61,w39_62,w39_63,w39_64,
		w39_65,w39_66,w39_67,w39_68,w39_69,w39_70,w39_71,w39_72,w39_73,w39_74,w39_75,w39_76,w39_77,w39_78,w39_79,w39_80,
		w39_81,w39_82,w39_83,w39_84,w39_85,w39_86,w39_87,w39_88,w39_89,w39_90,w39_91,w39_92,w39_93,w39_94,w39_95,w39_96,
		w39_97,w39_98,w39_99,w39_100,w39_101,w39_102,w39_103,w39_104,w39_105,w39_106,w39_107,w39_108,w39_109,w39_110,w39_111,w39_112,
		w39_113,w39_114,w39_115,w39_116,w39_117,w39_118,w39_119,w39_120,w39_121,w39_122,w39_123,w39_124,w39_125,w39_126,
	w40_0,w40_1,w40_2,w40_3,w40_4,w40_5,w40_6,w40_7,w40_8,w40_9,w40_10,w40_11,w40_12,w40_13,w40_14,w40_15,w40_16,
		w40_17,w40_18,w40_19,w40_20,w40_21,w40_22,w40_23,w40_24,w40_25,w40_26,w40_27,w40_28,w40_29,w40_30,w40_31,w40_32,
		w40_33,w40_34,w40_35,w40_36,w40_37,w40_38,w40_39,w40_40,w40_41,w40_42,w40_43,w40_44,w40_45,w40_46,w40_47,w40_48,
		w40_49,w40_50,w40_51,w40_52,w40_53,w40_54,w40_55,w40_56,w40_57,w40_58,w40_59,w40_60,w40_61,w40_62,w40_63,w40_64,
		w40_65,w40_66,w40_67,w40_68,w40_69,w40_70,w40_71,w40_72,w40_73,w40_74,w40_75,w40_76,w40_77,w40_78,w40_79,w40_80,
		w40_81,w40_82,w40_83,w40_84,w40_85,w40_86,w40_87,w40_88,w40_89,w40_90,w40_91,w40_92,w40_93,w40_94,w40_95,w40_96,
		w40_97,w40_98,w40_99,w40_100,w40_101,w40_102,w40_103,w40_104,w40_105,w40_106,w40_107,w40_108,w40_109,w40_110,w40_111,w40_112,
		w40_113,w40_114,w40_115,w40_116,w40_117,w40_118,w40_119,w40_120,w40_121,w40_122,w40_123,w40_124,w40_125,w40_126,
	w41_0,w41_1,w41_2,w41_3,w41_4,w41_5,w41_6,w41_7,w41_8,w41_9,w41_10,w41_11,w41_12,w41_13,w41_14,w41_15,w41_16,
		w41_17,w41_18,w41_19,w41_20,w41_21,w41_22,w41_23,w41_24,w41_25,w41_26,w41_27,w41_28,w41_29,w41_30,w41_31,w41_32,
		w41_33,w41_34,w41_35,w41_36,w41_37,w41_38,w41_39,w41_40,w41_41,w41_42,w41_43,w41_44,w41_45,w41_46,w41_47,w41_48,
		w41_49,w41_50,w41_51,w41_52,w41_53,w41_54,w41_55,w41_56,w41_57,w41_58,w41_59,w41_60,w41_61,w41_62,w41_63,w41_64,
		w41_65,w41_66,w41_67,w41_68,w41_69,w41_70,w41_71,w41_72,w41_73,w41_74,w41_75,w41_76,w41_77,w41_78,w41_79,w41_80,
		w41_81,w41_82,w41_83,w41_84,w41_85,w41_86,w41_87,w41_88,w41_89,w41_90,w41_91,w41_92,w41_93,w41_94,w41_95,w41_96,
		w41_97,w41_98,w41_99,w41_100,w41_101,w41_102,w41_103,w41_104,w41_105,w41_106,w41_107,w41_108,w41_109,w41_110,w41_111,w41_112,
		w41_113,w41_114,w41_115,w41_116,w41_117,w41_118,w41_119,w41_120,w41_121,w41_122,w41_123,w41_124,w41_125,w41_126,
	w42_0,w42_1,w42_2,w42_3,w42_4,w42_5,w42_6,w42_7,w42_8,w42_9,w42_10,w42_11,w42_12,w42_13,w42_14,w42_15,w42_16,
		w42_17,w42_18,w42_19,w42_20,w42_21,w42_22,w42_23,w42_24,w42_25,w42_26,w42_27,w42_28,w42_29,w42_30,w42_31,w42_32,
		w42_33,w42_34,w42_35,w42_36,w42_37,w42_38,w42_39,w42_40,w42_41,w42_42,w42_43,w42_44,w42_45,w42_46,w42_47,w42_48,
		w42_49,w42_50,w42_51,w42_52,w42_53,w42_54,w42_55,w42_56,w42_57,w42_58,w42_59,w42_60,w42_61,w42_62,w42_63,w42_64,
		w42_65,w42_66,w42_67,w42_68,w42_69,w42_70,w42_71,w42_72,w42_73,w42_74,w42_75,w42_76,w42_77,w42_78,w42_79,w42_80,
		w42_81,w42_82,w42_83,w42_84,w42_85,w42_86,w42_87,w42_88,w42_89,w42_90,w42_91,w42_92,w42_93,w42_94,w42_95,w42_96,
		w42_97,w42_98,w42_99,w42_100,w42_101,w42_102,w42_103,w42_104,w42_105,w42_106,w42_107,w42_108,w42_109,w42_110,w42_111,w42_112,
		w42_113,w42_114,w42_115,w42_116,w42_117,w42_118,w42_119,w42_120,w42_121,w42_122,w42_123,w42_124,w42_125,w42_126,
	w43_0,w43_1,w43_2,w43_3,w43_4,w43_5,w43_6,w43_7,w43_8,w43_9,w43_10,w43_11,w43_12,w43_13,w43_14,w43_15,w43_16,
		w43_17,w43_18,w43_19,w43_20,w43_21,w43_22,w43_23,w43_24,w43_25,w43_26,w43_27,w43_28,w43_29,w43_30,w43_31,w43_32,
		w43_33,w43_34,w43_35,w43_36,w43_37,w43_38,w43_39,w43_40,w43_41,w43_42,w43_43,w43_44,w43_45,w43_46,w43_47,w43_48,
		w43_49,w43_50,w43_51,w43_52,w43_53,w43_54,w43_55,w43_56,w43_57,w43_58,w43_59,w43_60,w43_61,w43_62,w43_63,w43_64,
		w43_65,w43_66,w43_67,w43_68,w43_69,w43_70,w43_71,w43_72,w43_73,w43_74,w43_75,w43_76,w43_77,w43_78,w43_79,w43_80,
		w43_81,w43_82,w43_83,w43_84,w43_85,w43_86,w43_87,w43_88,w43_89,w43_90,w43_91,w43_92,w43_93,w43_94,w43_95,w43_96,
		w43_97,w43_98,w43_99,w43_100,w43_101,w43_102,w43_103,w43_104,w43_105,w43_106,w43_107,w43_108,w43_109,w43_110,w43_111,w43_112,
		w43_113,w43_114,w43_115,w43_116,w43_117,w43_118,w43_119,w43_120,w43_121,w43_122,w43_123,w43_124,w43_125,w43_126,
	w44_0,w44_1,w44_2,w44_3,w44_4,w44_5,w44_6,w44_7,w44_8,w44_9,w44_10,w44_11,w44_12,w44_13,w44_14,w44_15,w44_16,
		w44_17,w44_18,w44_19,w44_20,w44_21,w44_22,w44_23,w44_24,w44_25,w44_26,w44_27,w44_28,w44_29,w44_30,w44_31,w44_32,
		w44_33,w44_34,w44_35,w44_36,w44_37,w44_38,w44_39,w44_40,w44_41,w44_42,w44_43,w44_44,w44_45,w44_46,w44_47,w44_48,
		w44_49,w44_50,w44_51,w44_52,w44_53,w44_54,w44_55,w44_56,w44_57,w44_58,w44_59,w44_60,w44_61,w44_62,w44_63,w44_64,
		w44_65,w44_66,w44_67,w44_68,w44_69,w44_70,w44_71,w44_72,w44_73,w44_74,w44_75,w44_76,w44_77,w44_78,w44_79,w44_80,
		w44_81,w44_82,w44_83,w44_84,w44_85,w44_86,w44_87,w44_88,w44_89,w44_90,w44_91,w44_92,w44_93,w44_94,w44_95,w44_96,
		w44_97,w44_98,w44_99,w44_100,w44_101,w44_102,w44_103,w44_104,w44_105,w44_106,w44_107,w44_108,w44_109,w44_110,w44_111,w44_112,
		w44_113,w44_114,w44_115,w44_116,w44_117,w44_118,w44_119,w44_120,w44_121,w44_122,w44_123,w44_124,w44_125,w44_126,
	w45_0,w45_1,w45_2,w45_3,w45_4,w45_5,w45_6,w45_7,w45_8,w45_9,w45_10,w45_11,w45_12,w45_13,w45_14,w45_15,w45_16,
		w45_17,w45_18,w45_19,w45_20,w45_21,w45_22,w45_23,w45_24,w45_25,w45_26,w45_27,w45_28,w45_29,w45_30,w45_31,w45_32,
		w45_33,w45_34,w45_35,w45_36,w45_37,w45_38,w45_39,w45_40,w45_41,w45_42,w45_43,w45_44,w45_45,w45_46,w45_47,w45_48,
		w45_49,w45_50,w45_51,w45_52,w45_53,w45_54,w45_55,w45_56,w45_57,w45_58,w45_59,w45_60,w45_61,w45_62,w45_63,w45_64,
		w45_65,w45_66,w45_67,w45_68,w45_69,w45_70,w45_71,w45_72,w45_73,w45_74,w45_75,w45_76,w45_77,w45_78,w45_79,w45_80,
		w45_81,w45_82,w45_83,w45_84,w45_85,w45_86,w45_87,w45_88,w45_89,w45_90,w45_91,w45_92,w45_93,w45_94,w45_95,w45_96,
		w45_97,w45_98,w45_99,w45_100,w45_101,w45_102,w45_103,w45_104,w45_105,w45_106,w45_107,w45_108,w45_109,w45_110,w45_111,w45_112,
		w45_113,w45_114,w45_115,w45_116,w45_117,w45_118,w45_119,w45_120,w45_121,w45_122,w45_123,w45_124,w45_125,w45_126,
	w46_0,w46_1,w46_2,w46_3,w46_4,w46_5,w46_6,w46_7,w46_8,w46_9,w46_10,w46_11,w46_12,w46_13,w46_14,w46_15,w46_16,
		w46_17,w46_18,w46_19,w46_20,w46_21,w46_22,w46_23,w46_24,w46_25,w46_26,w46_27,w46_28,w46_29,w46_30,w46_31,w46_32,
		w46_33,w46_34,w46_35,w46_36,w46_37,w46_38,w46_39,w46_40,w46_41,w46_42,w46_43,w46_44,w46_45,w46_46,w46_47,w46_48,
		w46_49,w46_50,w46_51,w46_52,w46_53,w46_54,w46_55,w46_56,w46_57,w46_58,w46_59,w46_60,w46_61,w46_62,w46_63,w46_64,
		w46_65,w46_66,w46_67,w46_68,w46_69,w46_70,w46_71,w46_72,w46_73,w46_74,w46_75,w46_76,w46_77,w46_78,w46_79,w46_80,
		w46_81,w46_82,w46_83,w46_84,w46_85,w46_86,w46_87,w46_88,w46_89,w46_90,w46_91,w46_92,w46_93,w46_94,w46_95,w46_96,
		w46_97,w46_98,w46_99,w46_100,w46_101,w46_102,w46_103,w46_104,w46_105,w46_106,w46_107,w46_108,w46_109,w46_110,w46_111,w46_112,
		w46_113,w46_114,w46_115,w46_116,w46_117,w46_118,w46_119,w46_120,w46_121,w46_122,w46_123,w46_124,w46_125,w46_126,
	w47_0,w47_1,w47_2,w47_3,w47_4,w47_5,w47_6,w47_7,w47_8,w47_9,w47_10,w47_11,w47_12,w47_13,w47_14,w47_15,w47_16,
		w47_17,w47_18,w47_19,w47_20,w47_21,w47_22,w47_23,w47_24,w47_25,w47_26,w47_27,w47_28,w47_29,w47_30,w47_31,w47_32,
		w47_33,w47_34,w47_35,w47_36,w47_37,w47_38,w47_39,w47_40,w47_41,w47_42,w47_43,w47_44,w47_45,w47_46,w47_47,w47_48,
		w47_49,w47_50,w47_51,w47_52,w47_53,w47_54,w47_55,w47_56,w47_57,w47_58,w47_59,w47_60,w47_61,w47_62,w47_63,w47_64,
		w47_65,w47_66,w47_67,w47_68,w47_69,w47_70,w47_71,w47_72,w47_73,w47_74,w47_75,w47_76,w47_77,w47_78,w47_79,w47_80,
		w47_81,w47_82,w47_83,w47_84,w47_85,w47_86,w47_87,w47_88,w47_89,w47_90,w47_91,w47_92,w47_93,w47_94,w47_95,w47_96,
		w47_97,w47_98,w47_99,w47_100,w47_101,w47_102,w47_103,w47_104,w47_105,w47_106,w47_107,w47_108,w47_109,w47_110,w47_111,w47_112,
		w47_113,w47_114,w47_115,w47_116,w47_117,w47_118,w47_119,w47_120,w47_121,w47_122,w47_123,w47_124,w47_125,w47_126,
	w48_0,w48_1,w48_2,w48_3,w48_4,w48_5,w48_6,w48_7,w48_8,w48_9,w48_10,w48_11,w48_12,w48_13,w48_14,w48_15,w48_16,
		w48_17,w48_18,w48_19,w48_20,w48_21,w48_22,w48_23,w48_24,w48_25,w48_26,w48_27,w48_28,w48_29,w48_30,w48_31,w48_32,
		w48_33,w48_34,w48_35,w48_36,w48_37,w48_38,w48_39,w48_40,w48_41,w48_42,w48_43,w48_44,w48_45,w48_46,w48_47,w48_48,
		w48_49,w48_50,w48_51,w48_52,w48_53,w48_54,w48_55,w48_56,w48_57,w48_58,w48_59,w48_60,w48_61,w48_62,w48_63,w48_64,
		w48_65,w48_66,w48_67,w48_68,w48_69,w48_70,w48_71,w48_72,w48_73,w48_74,w48_75,w48_76,w48_77,w48_78,w48_79,w48_80,
		w48_81,w48_82,w48_83,w48_84,w48_85,w48_86,w48_87,w48_88,w48_89,w48_90,w48_91,w48_92,w48_93,w48_94,w48_95,w48_96,
		w48_97,w48_98,w48_99,w48_100,w48_101,w48_102,w48_103,w48_104,w48_105,w48_106,w48_107,w48_108,w48_109,w48_110,w48_111,w48_112,
		w48_113,w48_114,w48_115,w48_116,w48_117,w48_118,w48_119,w48_120,w48_121,w48_122,w48_123,w48_124,w48_125,w48_126,
	w49_0,w49_1,w49_2,w49_3,w49_4,w49_5,w49_6,w49_7,w49_8,w49_9,w49_10,w49_11,w49_12,w49_13,w49_14,w49_15,w49_16,
		w49_17,w49_18,w49_19,w49_20,w49_21,w49_22,w49_23,w49_24,w49_25,w49_26,w49_27,w49_28,w49_29,w49_30,w49_31,w49_32,
		w49_33,w49_34,w49_35,w49_36,w49_37,w49_38,w49_39,w49_40,w49_41,w49_42,w49_43,w49_44,w49_45,w49_46,w49_47,w49_48,
		w49_49,w49_50,w49_51,w49_52,w49_53,w49_54,w49_55,w49_56,w49_57,w49_58,w49_59,w49_60,w49_61,w49_62,w49_63,w49_64,
		w49_65,w49_66,w49_67,w49_68,w49_69,w49_70,w49_71,w49_72,w49_73,w49_74,w49_75,w49_76,w49_77,w49_78,w49_79,w49_80,
		w49_81,w49_82,w49_83,w49_84,w49_85,w49_86,w49_87,w49_88,w49_89,w49_90,w49_91,w49_92,w49_93,w49_94,w49_95,w49_96,
		w49_97,w49_98,w49_99,w49_100,w49_101,w49_102,w49_103,w49_104,w49_105,w49_106,w49_107,w49_108,w49_109,w49_110,w49_111,w49_112,
		w49_113,w49_114,w49_115,w49_116,w49_117,w49_118,w49_119,w49_120,w49_121,w49_122,w49_123,w49_124,w49_125,w49_126,
	w50_0,w50_1,w50_2,w50_3,w50_4,w50_5,w50_6,w50_7,w50_8,w50_9,w50_10,w50_11,w50_12,w50_13,w50_14,w50_15,w50_16,
		w50_17,w50_18,w50_19,w50_20,w50_21,w50_22,w50_23,w50_24,w50_25,w50_26,w50_27,w50_28,w50_29,w50_30,w50_31,w50_32,
		w50_33,w50_34,w50_35,w50_36,w50_37,w50_38,w50_39,w50_40,w50_41,w50_42,w50_43,w50_44,w50_45,w50_46,w50_47,w50_48,
		w50_49,w50_50,w50_51,w50_52,w50_53,w50_54,w50_55,w50_56,w50_57,w50_58,w50_59,w50_60,w50_61,w50_62,w50_63,w50_64,
		w50_65,w50_66,w50_67,w50_68,w50_69,w50_70,w50_71,w50_72,w50_73,w50_74,w50_75,w50_76,w50_77,w50_78,w50_79,w50_80,
		w50_81,w50_82,w50_83,w50_84,w50_85,w50_86,w50_87,w50_88,w50_89,w50_90,w50_91,w50_92,w50_93,w50_94,w50_95,w50_96,
		w50_97,w50_98,w50_99,w50_100,w50_101,w50_102,w50_103,w50_104,w50_105,w50_106,w50_107,w50_108,w50_109,w50_110,w50_111,w50_112,
		w50_113,w50_114,w50_115,w50_116,w50_117,w50_118,w50_119,w50_120,w50_121,w50_122,w50_123,w50_124,w50_125,w50_126,
	w51_0,w51_1,w51_2,w51_3,w51_4,w51_5,w51_6,w51_7,w51_8,w51_9,w51_10,w51_11,w51_12,w51_13,w51_14,w51_15,w51_16,
		w51_17,w51_18,w51_19,w51_20,w51_21,w51_22,w51_23,w51_24,w51_25,w51_26,w51_27,w51_28,w51_29,w51_30,w51_31,w51_32,
		w51_33,w51_34,w51_35,w51_36,w51_37,w51_38,w51_39,w51_40,w51_41,w51_42,w51_43,w51_44,w51_45,w51_46,w51_47,w51_48,
		w51_49,w51_50,w51_51,w51_52,w51_53,w51_54,w51_55,w51_56,w51_57,w51_58,w51_59,w51_60,w51_61,w51_62,w51_63,w51_64,
		w51_65,w51_66,w51_67,w51_68,w51_69,w51_70,w51_71,w51_72,w51_73,w51_74,w51_75,w51_76,w51_77,w51_78,w51_79,w51_80,
		w51_81,w51_82,w51_83,w51_84,w51_85,w51_86,w51_87,w51_88,w51_89,w51_90,w51_91,w51_92,w51_93,w51_94,w51_95,w51_96,
		w51_97,w51_98,w51_99,w51_100,w51_101,w51_102,w51_103,w51_104,w51_105,w51_106,w51_107,w51_108,w51_109,w51_110,w51_111,w51_112,
		w51_113,w51_114,w51_115,w51_116,w51_117,w51_118,w51_119,w51_120,w51_121,w51_122,w51_123,w51_124,w51_125,w51_126,
	w52_0,w52_1,w52_2,w52_3,w52_4,w52_5,w52_6,w52_7,w52_8,w52_9,w52_10,w52_11,w52_12,w52_13,w52_14,w52_15,w52_16,
		w52_17,w52_18,w52_19,w52_20,w52_21,w52_22,w52_23,w52_24,w52_25,w52_26,w52_27,w52_28,w52_29,w52_30,w52_31,w52_32,
		w52_33,w52_34,w52_35,w52_36,w52_37,w52_38,w52_39,w52_40,w52_41,w52_42,w52_43,w52_44,w52_45,w52_46,w52_47,w52_48,
		w52_49,w52_50,w52_51,w52_52,w52_53,w52_54,w52_55,w52_56,w52_57,w52_58,w52_59,w52_60,w52_61,w52_62,w52_63,w52_64,
		w52_65,w52_66,w52_67,w52_68,w52_69,w52_70,w52_71,w52_72,w52_73,w52_74,w52_75,w52_76,w52_77,w52_78,w52_79,w52_80,
		w52_81,w52_82,w52_83,w52_84,w52_85,w52_86,w52_87,w52_88,w52_89,w52_90,w52_91,w52_92,w52_93,w52_94,w52_95,w52_96,
		w52_97,w52_98,w52_99,w52_100,w52_101,w52_102,w52_103,w52_104,w52_105,w52_106,w52_107,w52_108,w52_109,w52_110,w52_111,w52_112,
		w52_113,w52_114,w52_115,w52_116,w52_117,w52_118,w52_119,w52_120,w52_121,w52_122,w52_123,w52_124,w52_125,w52_126,
	w53_0,w53_1,w53_2,w53_3,w53_4,w53_5,w53_6,w53_7,w53_8,w53_9,w53_10,w53_11,w53_12,w53_13,w53_14,w53_15,w53_16,
		w53_17,w53_18,w53_19,w53_20,w53_21,w53_22,w53_23,w53_24,w53_25,w53_26,w53_27,w53_28,w53_29,w53_30,w53_31,w53_32,
		w53_33,w53_34,w53_35,w53_36,w53_37,w53_38,w53_39,w53_40,w53_41,w53_42,w53_43,w53_44,w53_45,w53_46,w53_47,w53_48,
		w53_49,w53_50,w53_51,w53_52,w53_53,w53_54,w53_55,w53_56,w53_57,w53_58,w53_59,w53_60,w53_61,w53_62,w53_63,w53_64,
		w53_65,w53_66,w53_67,w53_68,w53_69,w53_70,w53_71,w53_72,w53_73,w53_74,w53_75,w53_76,w53_77,w53_78,w53_79,w53_80,
		w53_81,w53_82,w53_83,w53_84,w53_85,w53_86,w53_87,w53_88,w53_89,w53_90,w53_91,w53_92,w53_93,w53_94,w53_95,w53_96,
		w53_97,w53_98,w53_99,w53_100,w53_101,w53_102,w53_103,w53_104,w53_105,w53_106,w53_107,w53_108,w53_109,w53_110,w53_111,w53_112,
		w53_113,w53_114,w53_115,w53_116,w53_117,w53_118,w53_119,w53_120,w53_121,w53_122,w53_123,w53_124,w53_125,w53_126,
	w54_0,w54_1,w54_2,w54_3,w54_4,w54_5,w54_6,w54_7,w54_8,w54_9,w54_10,w54_11,w54_12,w54_13,w54_14,w54_15,w54_16,
		w54_17,w54_18,w54_19,w54_20,w54_21,w54_22,w54_23,w54_24,w54_25,w54_26,w54_27,w54_28,w54_29,w54_30,w54_31,w54_32,
		w54_33,w54_34,w54_35,w54_36,w54_37,w54_38,w54_39,w54_40,w54_41,w54_42,w54_43,w54_44,w54_45,w54_46,w54_47,w54_48,
		w54_49,w54_50,w54_51,w54_52,w54_53,w54_54,w54_55,w54_56,w54_57,w54_58,w54_59,w54_60,w54_61,w54_62,w54_63,w54_64,
		w54_65,w54_66,w54_67,w54_68,w54_69,w54_70,w54_71,w54_72,w54_73,w54_74,w54_75,w54_76,w54_77,w54_78,w54_79,w54_80,
		w54_81,w54_82,w54_83,w54_84,w54_85,w54_86,w54_87,w54_88,w54_89,w54_90,w54_91,w54_92,w54_93,w54_94,w54_95,w54_96,
		w54_97,w54_98,w54_99,w54_100,w54_101,w54_102,w54_103,w54_104,w54_105,w54_106,w54_107,w54_108,w54_109,w54_110,w54_111,w54_112,
		w54_113,w54_114,w54_115,w54_116,w54_117,w54_118,w54_119,w54_120,w54_121,w54_122,w54_123,w54_124,w54_125,w54_126,
	w55_0,w55_1,w55_2,w55_3,w55_4,w55_5,w55_6,w55_7,w55_8,w55_9,w55_10,w55_11,w55_12,w55_13,w55_14,w55_15,w55_16,
		w55_17,w55_18,w55_19,w55_20,w55_21,w55_22,w55_23,w55_24,w55_25,w55_26,w55_27,w55_28,w55_29,w55_30,w55_31,w55_32,
		w55_33,w55_34,w55_35,w55_36,w55_37,w55_38,w55_39,w55_40,w55_41,w55_42,w55_43,w55_44,w55_45,w55_46,w55_47,w55_48,
		w55_49,w55_50,w55_51,w55_52,w55_53,w55_54,w55_55,w55_56,w55_57,w55_58,w55_59,w55_60,w55_61,w55_62,w55_63,w55_64,
		w55_65,w55_66,w55_67,w55_68,w55_69,w55_70,w55_71,w55_72,w55_73,w55_74,w55_75,w55_76,w55_77,w55_78,w55_79,w55_80,
		w55_81,w55_82,w55_83,w55_84,w55_85,w55_86,w55_87,w55_88,w55_89,w55_90,w55_91,w55_92,w55_93,w55_94,w55_95,w55_96,
		w55_97,w55_98,w55_99,w55_100,w55_101,w55_102,w55_103,w55_104,w55_105,w55_106,w55_107,w55_108,w55_109,w55_110,w55_111,w55_112,
		w55_113,w55_114,w55_115,w55_116,w55_117,w55_118,w55_119,w55_120,w55_121,w55_122,w55_123,w55_124,w55_125,w55_126,
	w56_0,w56_1,w56_2,w56_3,w56_4,w56_5,w56_6,w56_7,w56_8,w56_9,w56_10,w56_11,w56_12,w56_13,w56_14,w56_15,w56_16,
		w56_17,w56_18,w56_19,w56_20,w56_21,w56_22,w56_23,w56_24,w56_25,w56_26,w56_27,w56_28,w56_29,w56_30,w56_31,w56_32,
		w56_33,w56_34,w56_35,w56_36,w56_37,w56_38,w56_39,w56_40,w56_41,w56_42,w56_43,w56_44,w56_45,w56_46,w56_47,w56_48,
		w56_49,w56_50,w56_51,w56_52,w56_53,w56_54,w56_55,w56_56,w56_57,w56_58,w56_59,w56_60,w56_61,w56_62,w56_63,w56_64,
		w56_65,w56_66,w56_67,w56_68,w56_69,w56_70,w56_71,w56_72,w56_73,w56_74,w56_75,w56_76,w56_77,w56_78,w56_79,w56_80,
		w56_81,w56_82,w56_83,w56_84,w56_85,w56_86,w56_87,w56_88,w56_89,w56_90,w56_91,w56_92,w56_93,w56_94,w56_95,w56_96,
		w56_97,w56_98,w56_99,w56_100,w56_101,w56_102,w56_103,w56_104,w56_105,w56_106,w56_107,w56_108,w56_109,w56_110,w56_111,w56_112,
		w56_113,w56_114,w56_115,w56_116,w56_117,w56_118,w56_119,w56_120,w56_121,w56_122,w56_123,w56_124,w56_125,w56_126,
	w57_0,w57_1,w57_2,w57_3,w57_4,w57_5,w57_6,w57_7,w57_8,w57_9,w57_10,w57_11,w57_12,w57_13,w57_14,w57_15,w57_16,
		w57_17,w57_18,w57_19,w57_20,w57_21,w57_22,w57_23,w57_24,w57_25,w57_26,w57_27,w57_28,w57_29,w57_30,w57_31,w57_32,
		w57_33,w57_34,w57_35,w57_36,w57_37,w57_38,w57_39,w57_40,w57_41,w57_42,w57_43,w57_44,w57_45,w57_46,w57_47,w57_48,
		w57_49,w57_50,w57_51,w57_52,w57_53,w57_54,w57_55,w57_56,w57_57,w57_58,w57_59,w57_60,w57_61,w57_62,w57_63,w57_64,
		w57_65,w57_66,w57_67,w57_68,w57_69,w57_70,w57_71,w57_72,w57_73,w57_74,w57_75,w57_76,w57_77,w57_78,w57_79,w57_80,
		w57_81,w57_82,w57_83,w57_84,w57_85,w57_86,w57_87,w57_88,w57_89,w57_90,w57_91,w57_92,w57_93,w57_94,w57_95,w57_96,
		w57_97,w57_98,w57_99,w57_100,w57_101,w57_102,w57_103,w57_104,w57_105,w57_106,w57_107,w57_108,w57_109,w57_110,w57_111,w57_112,
		w57_113,w57_114,w57_115,w57_116,w57_117,w57_118,w57_119,w57_120,w57_121,w57_122,w57_123,w57_124,w57_125,w57_126,
	w58_0,w58_1,w58_2,w58_3,w58_4,w58_5,w58_6,w58_7,w58_8,w58_9,w58_10,w58_11,w58_12,w58_13,w58_14,w58_15,w58_16,
		w58_17,w58_18,w58_19,w58_20,w58_21,w58_22,w58_23,w58_24,w58_25,w58_26,w58_27,w58_28,w58_29,w58_30,w58_31,w58_32,
		w58_33,w58_34,w58_35,w58_36,w58_37,w58_38,w58_39,w58_40,w58_41,w58_42,w58_43,w58_44,w58_45,w58_46,w58_47,w58_48,
		w58_49,w58_50,w58_51,w58_52,w58_53,w58_54,w58_55,w58_56,w58_57,w58_58,w58_59,w58_60,w58_61,w58_62,w58_63,w58_64,
		w58_65,w58_66,w58_67,w58_68,w58_69,w58_70,w58_71,w58_72,w58_73,w58_74,w58_75,w58_76,w58_77,w58_78,w58_79,w58_80,
		w58_81,w58_82,w58_83,w58_84,w58_85,w58_86,w58_87,w58_88,w58_89,w58_90,w58_91,w58_92,w58_93,w58_94,w58_95,w58_96,
		w58_97,w58_98,w58_99,w58_100,w58_101,w58_102,w58_103,w58_104,w58_105,w58_106,w58_107,w58_108,w58_109,w58_110,w58_111,w58_112,
		w58_113,w58_114,w58_115,w58_116,w58_117,w58_118,w58_119,w58_120,w58_121,w58_122,w58_123,w58_124,w58_125,w58_126,
	w59_0,w59_1,w59_2,w59_3,w59_4,w59_5,w59_6,w59_7,w59_8,w59_9,w59_10,w59_11,w59_12,w59_13,w59_14,w59_15,w59_16,
		w59_17,w59_18,w59_19,w59_20,w59_21,w59_22,w59_23,w59_24,w59_25,w59_26,w59_27,w59_28,w59_29,w59_30,w59_31,w59_32,
		w59_33,w59_34,w59_35,w59_36,w59_37,w59_38,w59_39,w59_40,w59_41,w59_42,w59_43,w59_44,w59_45,w59_46,w59_47,w59_48,
		w59_49,w59_50,w59_51,w59_52,w59_53,w59_54,w59_55,w59_56,w59_57,w59_58,w59_59,w59_60,w59_61,w59_62,w59_63,w59_64,
		w59_65,w59_66,w59_67,w59_68,w59_69,w59_70,w59_71,w59_72,w59_73,w59_74,w59_75,w59_76,w59_77,w59_78,w59_79,w59_80,
		w59_81,w59_82,w59_83,w59_84,w59_85,w59_86,w59_87,w59_88,w59_89,w59_90,w59_91,w59_92,w59_93,w59_94,w59_95,w59_96,
		w59_97,w59_98,w59_99,w59_100,w59_101,w59_102,w59_103,w59_104,w59_105,w59_106,w59_107,w59_108,w59_109,w59_110,w59_111,w59_112,
		w59_113,w59_114,w59_115,w59_116,w59_117,w59_118,w59_119,w59_120,w59_121,w59_122,w59_123,w59_124,w59_125,w59_126,
	w60_0,w60_1,w60_2,w60_3,w60_4,w60_5,w60_6,w60_7,w60_8,w60_9,w60_10,w60_11,w60_12,w60_13,w60_14,w60_15,w60_16,
		w60_17,w60_18,w60_19,w60_20,w60_21,w60_22,w60_23,w60_24,w60_25,w60_26,w60_27,w60_28,w60_29,w60_30,w60_31,w60_32,
		w60_33,w60_34,w60_35,w60_36,w60_37,w60_38,w60_39,w60_40,w60_41,w60_42,w60_43,w60_44,w60_45,w60_46,w60_47,w60_48,
		w60_49,w60_50,w60_51,w60_52,w60_53,w60_54,w60_55,w60_56,w60_57,w60_58,w60_59,w60_60,w60_61,w60_62,w60_63,w60_64,
		w60_65,w60_66,w60_67,w60_68,w60_69,w60_70,w60_71,w60_72,w60_73,w60_74,w60_75,w60_76,w60_77,w60_78,w60_79,w60_80,
		w60_81,w60_82,w60_83,w60_84,w60_85,w60_86,w60_87,w60_88,w60_89,w60_90,w60_91,w60_92,w60_93,w60_94,w60_95,w60_96,
		w60_97,w60_98,w60_99,w60_100,w60_101,w60_102,w60_103,w60_104,w60_105,w60_106,w60_107,w60_108,w60_109,w60_110,w60_111,w60_112,
		w60_113,w60_114,w60_115,w60_116,w60_117,w60_118,w60_119,w60_120,w60_121,w60_122,w60_123,w60_124,w60_125,w60_126,
	w61_0,w61_1,w61_2,w61_3,w61_4,w61_5,w61_6,w61_7,w61_8,w61_9,w61_10,w61_11,w61_12,w61_13,w61_14,w61_15,w61_16,
		w61_17,w61_18,w61_19,w61_20,w61_21,w61_22,w61_23,w61_24,w61_25,w61_26,w61_27,w61_28,w61_29,w61_30,w61_31,w61_32,
		w61_33,w61_34,w61_35,w61_36,w61_37,w61_38,w61_39,w61_40,w61_41,w61_42,w61_43,w61_44,w61_45,w61_46,w61_47,w61_48,
		w61_49,w61_50,w61_51,w61_52,w61_53,w61_54,w61_55,w61_56,w61_57,w61_58,w61_59,w61_60,w61_61,w61_62,w61_63,w61_64,
		w61_65,w61_66,w61_67,w61_68,w61_69,w61_70,w61_71,w61_72,w61_73,w61_74,w61_75,w61_76,w61_77,w61_78,w61_79,w61_80,
		w61_81,w61_82,w61_83,w61_84,w61_85,w61_86,w61_87,w61_88,w61_89,w61_90,w61_91,w61_92,w61_93,w61_94,w61_95,w61_96,
		w61_97,w61_98,w61_99,w61_100,w61_101,w61_102,w61_103,w61_104,w61_105,w61_106,w61_107,w61_108,w61_109,w61_110,w61_111,w61_112,
		w61_113,w61_114,w61_115,w61_116,w61_117,w61_118,w61_119,w61_120,w61_121,w61_122,w61_123,w61_124,w61_125,w61_126,
	w62_0,w62_1,w62_2,w62_3,w62_4,w62_5,w62_6,w62_7,w62_8,w62_9,w62_10,w62_11,w62_12,w62_13,w62_14,w62_15,w62_16,
		w62_17,w62_18,w62_19,w62_20,w62_21,w62_22,w62_23,w62_24,w62_25,w62_26,w62_27,w62_28,w62_29,w62_30,w62_31,w62_32,
		w62_33,w62_34,w62_35,w62_36,w62_37,w62_38,w62_39,w62_40,w62_41,w62_42,w62_43,w62_44,w62_45,w62_46,w62_47,w62_48,
		w62_49,w62_50,w62_51,w62_52,w62_53,w62_54,w62_55,w62_56,w62_57,w62_58,w62_59,w62_60,w62_61,w62_62,w62_63,w62_64,
		w62_65,w62_66,w62_67,w62_68,w62_69,w62_70,w62_71,w62_72,w62_73,w62_74,w62_75,w62_76,w62_77,w62_78,w62_79,w62_80,
		w62_81,w62_82,w62_83,w62_84,w62_85,w62_86,w62_87,w62_88,w62_89,w62_90,w62_91,w62_92,w62_93,w62_94,w62_95,w62_96,
		w62_97,w62_98,w62_99,w62_100,w62_101,w62_102,w62_103,w62_104,w62_105,w62_106,w62_107,w62_108,w62_109,w62_110,w62_111,w62_112,
		w62_113,w62_114,w62_115,w62_116,w62_117,w62_118,w62_119,w62_120,w62_121,w62_122,w62_123,w62_124,w62_125,w62_126,
	w63_0,w63_1,w63_2,w63_3,w63_4,w63_5,w63_6,w63_7,w63_8,w63_9,w63_10,w63_11,w63_12,w63_13,w63_14,w63_15,w63_16,
		w63_17,w63_18,w63_19,w63_20,w63_21,w63_22,w63_23,w63_24,w63_25,w63_26,w63_27,w63_28,w63_29,w63_30,w63_31,w63_32,
		w63_33,w63_34,w63_35,w63_36,w63_37,w63_38,w63_39,w63_40,w63_41,w63_42,w63_43,w63_44,w63_45,w63_46,w63_47,w63_48,
		w63_49,w63_50,w63_51,w63_52,w63_53,w63_54,w63_55,w63_56,w63_57,w63_58,w63_59,w63_60,w63_61,w63_62,w63_63,w63_64,
		w63_65,w63_66,w63_67,w63_68,w63_69,w63_70,w63_71,w63_72,w63_73,w63_74,w63_75,w63_76,w63_77,w63_78,w63_79,w63_80,
		w63_81,w63_82,w63_83,w63_84,w63_85,w63_86,w63_87,w63_88,w63_89,w63_90,w63_91,w63_92,w63_93,w63_94,w63_95,w63_96,
		w63_97,w63_98,w63_99,w63_100,w63_101,w63_102,w63_103,w63_104,w63_105,w63_106,w63_107,w63_108,w63_109,w63_110,w63_111,w63_112,
		w63_113,w63_114,w63_115,w63_116,w63_117,w63_118,w63_119,w63_120,w63_121,w63_122,w63_123,w63_124,w63_125,w63_126,
	w64_0,w64_1,w64_2,w64_3,w64_4,w64_5,w64_6,w64_7,w64_8,w64_9,w64_10,w64_11,w64_12,w64_13,w64_14,w64_15,w64_16,
		w64_17,w64_18,w64_19,w64_20,w64_21,w64_22,w64_23,w64_24,w64_25,w64_26,w64_27,w64_28,w64_29,w64_30,w64_31,w64_32,
		w64_33,w64_34,w64_35,w64_36,w64_37,w64_38,w64_39,w64_40,w64_41,w64_42,w64_43,w64_44,w64_45,w64_46,w64_47,w64_48,
		w64_49,w64_50,w64_51,w64_52,w64_53,w64_54,w64_55,w64_56,w64_57,w64_58,w64_59,w64_60,w64_61,w64_62,w64_63,w64_64,
		w64_65,w64_66,w64_67,w64_68,w64_69,w64_70,w64_71,w64_72,w64_73,w64_74,w64_75,w64_76,w64_77,w64_78,w64_79,w64_80,
		w64_81,w64_82,w64_83,w64_84,w64_85,w64_86,w64_87,w64_88,w64_89,w64_90,w64_91,w64_92,w64_93,w64_94,w64_95,w64_96,
		w64_97,w64_98,w64_99,w64_100,w64_101,w64_102,w64_103,w64_104,w64_105,w64_106,w64_107,w64_108,w64_109,w64_110,w64_111,w64_112,
		w64_113,w64_114,w64_115,w64_116,w64_117,w64_118,w64_119,w64_120,w64_121,w64_122,w64_123,w64_124,w64_125,w64_126,
	w65_0,w65_1,w65_2,w65_3,w65_4,w65_5,w65_6,w65_7,w65_8,w65_9,w65_10,w65_11,w65_12,w65_13,w65_14,w65_15,w65_16,
		w65_17,w65_18,w65_19,w65_20,w65_21,w65_22,w65_23,w65_24,w65_25,w65_26,w65_27,w65_28,w65_29,w65_30,w65_31,w65_32,
		w65_33,w65_34,w65_35,w65_36,w65_37,w65_38,w65_39,w65_40,w65_41,w65_42,w65_43,w65_44,w65_45,w65_46,w65_47,w65_48,
		w65_49,w65_50,w65_51,w65_52,w65_53,w65_54,w65_55,w65_56,w65_57,w65_58,w65_59,w65_60,w65_61,w65_62,w65_63,w65_64,
		w65_65,w65_66,w65_67,w65_68,w65_69,w65_70,w65_71,w65_72,w65_73,w65_74,w65_75,w65_76,w65_77,w65_78,w65_79,w65_80,
		w65_81,w65_82,w65_83,w65_84,w65_85,w65_86,w65_87,w65_88,w65_89,w65_90,w65_91,w65_92,w65_93,w65_94,w65_95,w65_96,
		w65_97,w65_98,w65_99,w65_100,w65_101,w65_102,w65_103,w65_104,w65_105,w65_106,w65_107,w65_108,w65_109,w65_110,w65_111,w65_112,
		w65_113,w65_114,w65_115,w65_116,w65_117,w65_118,w65_119,w65_120,w65_121,w65_122,w65_123,w65_124,w65_125,w65_126,
	w66_0,w66_1,w66_2,w66_3,w66_4,w66_5,w66_6,w66_7,w66_8,w66_9,w66_10,w66_11,w66_12,w66_13,w66_14,w66_15,w66_16,
		w66_17,w66_18,w66_19,w66_20,w66_21,w66_22,w66_23,w66_24,w66_25,w66_26,w66_27,w66_28,w66_29,w66_30,w66_31,w66_32,
		w66_33,w66_34,w66_35,w66_36,w66_37,w66_38,w66_39,w66_40,w66_41,w66_42,w66_43,w66_44,w66_45,w66_46,w66_47,w66_48,
		w66_49,w66_50,w66_51,w66_52,w66_53,w66_54,w66_55,w66_56,w66_57,w66_58,w66_59,w66_60,w66_61,w66_62,w66_63,w66_64,
		w66_65,w66_66,w66_67,w66_68,w66_69,w66_70,w66_71,w66_72,w66_73,w66_74,w66_75,w66_76,w66_77,w66_78,w66_79,w66_80,
		w66_81,w66_82,w66_83,w66_84,w66_85,w66_86,w66_87,w66_88,w66_89,w66_90,w66_91,w66_92,w66_93,w66_94,w66_95,w66_96,
		w66_97,w66_98,w66_99,w66_100,w66_101,w66_102,w66_103,w66_104,w66_105,w66_106,w66_107,w66_108,w66_109,w66_110,w66_111,w66_112,
		w66_113,w66_114,w66_115,w66_116,w66_117,w66_118,w66_119,w66_120,w66_121,w66_122,w66_123,w66_124,w66_125,w66_126,
	w67_0,w67_1,w67_2,w67_3,w67_4,w67_5,w67_6,w67_7,w67_8,w67_9,w67_10,w67_11,w67_12,w67_13,w67_14,w67_15,w67_16,
		w67_17,w67_18,w67_19,w67_20,w67_21,w67_22,w67_23,w67_24,w67_25,w67_26,w67_27,w67_28,w67_29,w67_30,w67_31,w67_32,
		w67_33,w67_34,w67_35,w67_36,w67_37,w67_38,w67_39,w67_40,w67_41,w67_42,w67_43,w67_44,w67_45,w67_46,w67_47,w67_48,
		w67_49,w67_50,w67_51,w67_52,w67_53,w67_54,w67_55,w67_56,w67_57,w67_58,w67_59,w67_60,w67_61,w67_62,w67_63,w67_64,
		w67_65,w67_66,w67_67,w67_68,w67_69,w67_70,w67_71,w67_72,w67_73,w67_74,w67_75,w67_76,w67_77,w67_78,w67_79,w67_80,
		w67_81,w67_82,w67_83,w67_84,w67_85,w67_86,w67_87,w67_88,w67_89,w67_90,w67_91,w67_92,w67_93,w67_94,w67_95,w67_96,
		w67_97,w67_98,w67_99,w67_100,w67_101,w67_102,w67_103,w67_104,w67_105,w67_106,w67_107,w67_108,w67_109,w67_110,w67_111,w67_112,
		w67_113,w67_114,w67_115,w67_116,w67_117,w67_118,w67_119,w67_120,w67_121,w67_122,w67_123,w67_124,w67_125,w67_126,
	w68_0,w68_1,w68_2,w68_3,w68_4,w68_5,w68_6,w68_7,w68_8,w68_9,w68_10,w68_11,w68_12,w68_13,w68_14,w68_15,w68_16,
		w68_17,w68_18,w68_19,w68_20,w68_21,w68_22,w68_23,w68_24,w68_25,w68_26,w68_27,w68_28,w68_29,w68_30,w68_31,w68_32,
		w68_33,w68_34,w68_35,w68_36,w68_37,w68_38,w68_39,w68_40,w68_41,w68_42,w68_43,w68_44,w68_45,w68_46,w68_47,w68_48,
		w68_49,w68_50,w68_51,w68_52,w68_53,w68_54,w68_55,w68_56,w68_57,w68_58,w68_59,w68_60,w68_61,w68_62,w68_63,w68_64,
		w68_65,w68_66,w68_67,w68_68,w68_69,w68_70,w68_71,w68_72,w68_73,w68_74,w68_75,w68_76,w68_77,w68_78,w68_79,w68_80,
		w68_81,w68_82,w68_83,w68_84,w68_85,w68_86,w68_87,w68_88,w68_89,w68_90,w68_91,w68_92,w68_93,w68_94,w68_95,w68_96,
		w68_97,w68_98,w68_99,w68_100,w68_101,w68_102,w68_103,w68_104,w68_105,w68_106,w68_107,w68_108,w68_109,w68_110,w68_111,w68_112,
		w68_113,w68_114,w68_115,w68_116,w68_117,w68_118,w68_119,w68_120,w68_121,w68_122,w68_123,w68_124,w68_125,w68_126,
	w69_0,w69_1,w69_2,w69_3,w69_4,w69_5,w69_6,w69_7,w69_8,w69_9,w69_10,w69_11,w69_12,w69_13,w69_14,w69_15,w69_16,
		w69_17,w69_18,w69_19,w69_20,w69_21,w69_22,w69_23,w69_24,w69_25,w69_26,w69_27,w69_28,w69_29,w69_30,w69_31,w69_32,
		w69_33,w69_34,w69_35,w69_36,w69_37,w69_38,w69_39,w69_40,w69_41,w69_42,w69_43,w69_44,w69_45,w69_46,w69_47,w69_48,
		w69_49,w69_50,w69_51,w69_52,w69_53,w69_54,w69_55,w69_56,w69_57,w69_58,w69_59,w69_60,w69_61,w69_62,w69_63,w69_64,
		w69_65,w69_66,w69_67,w69_68,w69_69,w69_70,w69_71,w69_72,w69_73,w69_74,w69_75,w69_76,w69_77,w69_78,w69_79,w69_80,
		w69_81,w69_82,w69_83,w69_84,w69_85,w69_86,w69_87,w69_88,w69_89,w69_90,w69_91,w69_92,w69_93,w69_94,w69_95,w69_96,
		w69_97,w69_98,w69_99,w69_100,w69_101,w69_102,w69_103,w69_104,w69_105,w69_106,w69_107,w69_108,w69_109,w69_110,w69_111,w69_112,
		w69_113,w69_114,w69_115,w69_116,w69_117,w69_118,w69_119,w69_120,w69_121,w69_122,w69_123,w69_124,w69_125,w69_126,
	w70_0,w70_1,w70_2,w70_3,w70_4,w70_5,w70_6,w70_7,w70_8,w70_9,w70_10,w70_11,w70_12,w70_13,w70_14,w70_15,w70_16,
		w70_17,w70_18,w70_19,w70_20,w70_21,w70_22,w70_23,w70_24,w70_25,w70_26,w70_27,w70_28,w70_29,w70_30,w70_31,w70_32,
		w70_33,w70_34,w70_35,w70_36,w70_37,w70_38,w70_39,w70_40,w70_41,w70_42,w70_43,w70_44,w70_45,w70_46,w70_47,w70_48,
		w70_49,w70_50,w70_51,w70_52,w70_53,w70_54,w70_55,w70_56,w70_57,w70_58,w70_59,w70_60,w70_61,w70_62,w70_63,w70_64,
		w70_65,w70_66,w70_67,w70_68,w70_69,w70_70,w70_71,w70_72,w70_73,w70_74,w70_75,w70_76,w70_77,w70_78,w70_79,w70_80,
		w70_81,w70_82,w70_83,w70_84,w70_85,w70_86,w70_87,w70_88,w70_89,w70_90,w70_91,w70_92,w70_93,w70_94,w70_95,w70_96,
		w70_97,w70_98,w70_99,w70_100,w70_101,w70_102,w70_103,w70_104,w70_105,w70_106,w70_107,w70_108,w70_109,w70_110,w70_111,w70_112,
		w70_113,w70_114,w70_115,w70_116,w70_117,w70_118,w70_119,w70_120,w70_121,w70_122,w70_123,w70_124,w70_125,w70_126,
	w71_0,w71_1,w71_2,w71_3,w71_4,w71_5,w71_6,w71_7,w71_8,w71_9,w71_10,w71_11,w71_12,w71_13,w71_14,w71_15,w71_16,
		w71_17,w71_18,w71_19,w71_20,w71_21,w71_22,w71_23,w71_24,w71_25,w71_26,w71_27,w71_28,w71_29,w71_30,w71_31,w71_32,
		w71_33,w71_34,w71_35,w71_36,w71_37,w71_38,w71_39,w71_40,w71_41,w71_42,w71_43,w71_44,w71_45,w71_46,w71_47,w71_48,
		w71_49,w71_50,w71_51,w71_52,w71_53,w71_54,w71_55,w71_56,w71_57,w71_58,w71_59,w71_60,w71_61,w71_62,w71_63,w71_64,
		w71_65,w71_66,w71_67,w71_68,w71_69,w71_70,w71_71,w71_72,w71_73,w71_74,w71_75,w71_76,w71_77,w71_78,w71_79,w71_80,
		w71_81,w71_82,w71_83,w71_84,w71_85,w71_86,w71_87,w71_88,w71_89,w71_90,w71_91,w71_92,w71_93,w71_94,w71_95,w71_96,
		w71_97,w71_98,w71_99,w71_100,w71_101,w71_102,w71_103,w71_104,w71_105,w71_106,w71_107,w71_108,w71_109,w71_110,w71_111,w71_112,
		w71_113,w71_114,w71_115,w71_116,w71_117,w71_118,w71_119,w71_120,w71_121,w71_122,w71_123,w71_124,w71_125,w71_126,
	w72_0,w72_1,w72_2,w72_3,w72_4,w72_5,w72_6,w72_7,w72_8,w72_9,w72_10,w72_11,w72_12,w72_13,w72_14,w72_15,w72_16,
		w72_17,w72_18,w72_19,w72_20,w72_21,w72_22,w72_23,w72_24,w72_25,w72_26,w72_27,w72_28,w72_29,w72_30,w72_31,w72_32,
		w72_33,w72_34,w72_35,w72_36,w72_37,w72_38,w72_39,w72_40,w72_41,w72_42,w72_43,w72_44,w72_45,w72_46,w72_47,w72_48,
		w72_49,w72_50,w72_51,w72_52,w72_53,w72_54,w72_55,w72_56,w72_57,w72_58,w72_59,w72_60,w72_61,w72_62,w72_63,w72_64,
		w72_65,w72_66,w72_67,w72_68,w72_69,w72_70,w72_71,w72_72,w72_73,w72_74,w72_75,w72_76,w72_77,w72_78,w72_79,w72_80,
		w72_81,w72_82,w72_83,w72_84,w72_85,w72_86,w72_87,w72_88,w72_89,w72_90,w72_91,w72_92,w72_93,w72_94,w72_95,w72_96,
		w72_97,w72_98,w72_99,w72_100,w72_101,w72_102,w72_103,w72_104,w72_105,w72_106,w72_107,w72_108,w72_109,w72_110,w72_111,w72_112,
		w72_113,w72_114,w72_115,w72_116,w72_117,w72_118,w72_119,w72_120,w72_121,w72_122,w72_123,w72_124,w72_125,w72_126,
	w73_0,w73_1,w73_2,w73_3,w73_4,w73_5,w73_6,w73_7,w73_8,w73_9,w73_10,w73_11,w73_12,w73_13,w73_14,w73_15,w73_16,
		w73_17,w73_18,w73_19,w73_20,w73_21,w73_22,w73_23,w73_24,w73_25,w73_26,w73_27,w73_28,w73_29,w73_30,w73_31,w73_32,
		w73_33,w73_34,w73_35,w73_36,w73_37,w73_38,w73_39,w73_40,w73_41,w73_42,w73_43,w73_44,w73_45,w73_46,w73_47,w73_48,
		w73_49,w73_50,w73_51,w73_52,w73_53,w73_54,w73_55,w73_56,w73_57,w73_58,w73_59,w73_60,w73_61,w73_62,w73_63,w73_64,
		w73_65,w73_66,w73_67,w73_68,w73_69,w73_70,w73_71,w73_72,w73_73,w73_74,w73_75,w73_76,w73_77,w73_78,w73_79,w73_80,
		w73_81,w73_82,w73_83,w73_84,w73_85,w73_86,w73_87,w73_88,w73_89,w73_90,w73_91,w73_92,w73_93,w73_94,w73_95,w73_96,
		w73_97,w73_98,w73_99,w73_100,w73_101,w73_102,w73_103,w73_104,w73_105,w73_106,w73_107,w73_108,w73_109,w73_110,w73_111,w73_112,
		w73_113,w73_114,w73_115,w73_116,w73_117,w73_118,w73_119,w73_120,w73_121,w73_122,w73_123,w73_124,w73_125,w73_126,
	w74_0,w74_1,w74_2,w74_3,w74_4,w74_5,w74_6,w74_7,w74_8,w74_9,w74_10,w74_11,w74_12,w74_13,w74_14,w74_15,w74_16,
		w74_17,w74_18,w74_19,w74_20,w74_21,w74_22,w74_23,w74_24,w74_25,w74_26,w74_27,w74_28,w74_29,w74_30,w74_31,w74_32,
		w74_33,w74_34,w74_35,w74_36,w74_37,w74_38,w74_39,w74_40,w74_41,w74_42,w74_43,w74_44,w74_45,w74_46,w74_47,w74_48,
		w74_49,w74_50,w74_51,w74_52,w74_53,w74_54,w74_55,w74_56,w74_57,w74_58,w74_59,w74_60,w74_61,w74_62,w74_63,w74_64,
		w74_65,w74_66,w74_67,w74_68,w74_69,w74_70,w74_71,w74_72,w74_73,w74_74,w74_75,w74_76,w74_77,w74_78,w74_79,w74_80,
		w74_81,w74_82,w74_83,w74_84,w74_85,w74_86,w74_87,w74_88,w74_89,w74_90,w74_91,w74_92,w74_93,w74_94,w74_95,w74_96,
		w74_97,w74_98,w74_99,w74_100,w74_101,w74_102,w74_103,w74_104,w74_105,w74_106,w74_107,w74_108,w74_109,w74_110,w74_111,w74_112,
		w74_113,w74_114,w74_115,w74_116,w74_117,w74_118,w74_119,w74_120,w74_121,w74_122,w74_123,w74_124,w74_125,w74_126,
	w75_0,w75_1,w75_2,w75_3,w75_4,w75_5,w75_6,w75_7,w75_8,w75_9,w75_10,w75_11,w75_12,w75_13,w75_14,w75_15,w75_16,
		w75_17,w75_18,w75_19,w75_20,w75_21,w75_22,w75_23,w75_24,w75_25,w75_26,w75_27,w75_28,w75_29,w75_30,w75_31,w75_32,
		w75_33,w75_34,w75_35,w75_36,w75_37,w75_38,w75_39,w75_40,w75_41,w75_42,w75_43,w75_44,w75_45,w75_46,w75_47,w75_48,
		w75_49,w75_50,w75_51,w75_52,w75_53,w75_54,w75_55,w75_56,w75_57,w75_58,w75_59,w75_60,w75_61,w75_62,w75_63,w75_64,
		w75_65,w75_66,w75_67,w75_68,w75_69,w75_70,w75_71,w75_72,w75_73,w75_74,w75_75,w75_76,w75_77,w75_78,w75_79,w75_80,
		w75_81,w75_82,w75_83,w75_84,w75_85,w75_86,w75_87,w75_88,w75_89,w75_90,w75_91,w75_92,w75_93,w75_94,w75_95,w75_96,
		w75_97,w75_98,w75_99,w75_100,w75_101,w75_102,w75_103,w75_104,w75_105,w75_106,w75_107,w75_108,w75_109,w75_110,w75_111,w75_112,
		w75_113,w75_114,w75_115,w75_116,w75_117,w75_118,w75_119,w75_120,w75_121,w75_122,w75_123,w75_124,w75_125,w75_126,
	w76_0,w76_1,w76_2,w76_3,w76_4,w76_5,w76_6,w76_7,w76_8,w76_9,w76_10,w76_11,w76_12,w76_13,w76_14,w76_15,w76_16,
		w76_17,w76_18,w76_19,w76_20,w76_21,w76_22,w76_23,w76_24,w76_25,w76_26,w76_27,w76_28,w76_29,w76_30,w76_31,w76_32,
		w76_33,w76_34,w76_35,w76_36,w76_37,w76_38,w76_39,w76_40,w76_41,w76_42,w76_43,w76_44,w76_45,w76_46,w76_47,w76_48,
		w76_49,w76_50,w76_51,w76_52,w76_53,w76_54,w76_55,w76_56,w76_57,w76_58,w76_59,w76_60,w76_61,w76_62,w76_63,w76_64,
		w76_65,w76_66,w76_67,w76_68,w76_69,w76_70,w76_71,w76_72,w76_73,w76_74,w76_75,w76_76,w76_77,w76_78,w76_79,w76_80,
		w76_81,w76_82,w76_83,w76_84,w76_85,w76_86,w76_87,w76_88,w76_89,w76_90,w76_91,w76_92,w76_93,w76_94,w76_95,w76_96,
		w76_97,w76_98,w76_99,w76_100,w76_101,w76_102,w76_103,w76_104,w76_105,w76_106,w76_107,w76_108,w76_109,w76_110,w76_111,w76_112,
		w76_113,w76_114,w76_115,w76_116,w76_117,w76_118,w76_119,w76_120,w76_121,w76_122,w76_123,w76_124,w76_125,w76_126,
	w77_0,w77_1,w77_2,w77_3,w77_4,w77_5,w77_6,w77_7,w77_8,w77_9,w77_10,w77_11,w77_12,w77_13,w77_14,w77_15,w77_16,
		w77_17,w77_18,w77_19,w77_20,w77_21,w77_22,w77_23,w77_24,w77_25,w77_26,w77_27,w77_28,w77_29,w77_30,w77_31,w77_32,
		w77_33,w77_34,w77_35,w77_36,w77_37,w77_38,w77_39,w77_40,w77_41,w77_42,w77_43,w77_44,w77_45,w77_46,w77_47,w77_48,
		w77_49,w77_50,w77_51,w77_52,w77_53,w77_54,w77_55,w77_56,w77_57,w77_58,w77_59,w77_60,w77_61,w77_62,w77_63,w77_64,
		w77_65,w77_66,w77_67,w77_68,w77_69,w77_70,w77_71,w77_72,w77_73,w77_74,w77_75,w77_76,w77_77,w77_78,w77_79,w77_80,
		w77_81,w77_82,w77_83,w77_84,w77_85,w77_86,w77_87,w77_88,w77_89,w77_90,w77_91,w77_92,w77_93,w77_94,w77_95,w77_96,
		w77_97,w77_98,w77_99,w77_100,w77_101,w77_102,w77_103,w77_104,w77_105,w77_106,w77_107,w77_108,w77_109,w77_110,w77_111,w77_112,
		w77_113,w77_114,w77_115,w77_116,w77_117,w77_118,w77_119,w77_120,w77_121,w77_122,w77_123,w77_124,w77_125,w77_126,
	w78_0,w78_1,w78_2,w78_3,w78_4,w78_5,w78_6,w78_7,w78_8,w78_9,w78_10,w78_11,w78_12,w78_13,w78_14,w78_15,w78_16,
		w78_17,w78_18,w78_19,w78_20,w78_21,w78_22,w78_23,w78_24,w78_25,w78_26,w78_27,w78_28,w78_29,w78_30,w78_31,w78_32,
		w78_33,w78_34,w78_35,w78_36,w78_37,w78_38,w78_39,w78_40,w78_41,w78_42,w78_43,w78_44,w78_45,w78_46,w78_47,w78_48,
		w78_49,w78_50,w78_51,w78_52,w78_53,w78_54,w78_55,w78_56,w78_57,w78_58,w78_59,w78_60,w78_61,w78_62,w78_63,w78_64,
		w78_65,w78_66,w78_67,w78_68,w78_69,w78_70,w78_71,w78_72,w78_73,w78_74,w78_75,w78_76,w78_77,w78_78,w78_79,w78_80,
		w78_81,w78_82,w78_83,w78_84,w78_85,w78_86,w78_87,w78_88,w78_89,w78_90,w78_91,w78_92,w78_93,w78_94,w78_95,w78_96,
		w78_97,w78_98,w78_99,w78_100,w78_101,w78_102,w78_103,w78_104,w78_105,w78_106,w78_107,w78_108,w78_109,w78_110,w78_111,w78_112,
		w78_113,w78_114,w78_115,w78_116,w78_117,w78_118,w78_119,w78_120,w78_121,w78_122,w78_123,w78_124,w78_125,w78_126,
	w79_0,w79_1,w79_2,w79_3,w79_4,w79_5,w79_6,w79_7,w79_8,w79_9,w79_10,w79_11,w79_12,w79_13,w79_14,w79_15,w79_16,
		w79_17,w79_18,w79_19,w79_20,w79_21,w79_22,w79_23,w79_24,w79_25,w79_26,w79_27,w79_28,w79_29,w79_30,w79_31,w79_32,
		w79_33,w79_34,w79_35,w79_36,w79_37,w79_38,w79_39,w79_40,w79_41,w79_42,w79_43,w79_44,w79_45,w79_46,w79_47,w79_48,
		w79_49,w79_50,w79_51,w79_52,w79_53,w79_54,w79_55,w79_56,w79_57,w79_58,w79_59,w79_60,w79_61,w79_62,w79_63,w79_64,
		w79_65,w79_66,w79_67,w79_68,w79_69,w79_70,w79_71,w79_72,w79_73,w79_74,w79_75,w79_76,w79_77,w79_78,w79_79,w79_80,
		w79_81,w79_82,w79_83,w79_84,w79_85,w79_86,w79_87,w79_88,w79_89,w79_90,w79_91,w79_92,w79_93,w79_94,w79_95,w79_96,
		w79_97,w79_98,w79_99,w79_100,w79_101,w79_102,w79_103,w79_104,w79_105,w79_106,w79_107,w79_108,w79_109,w79_110,w79_111,w79_112,
		w79_113,w79_114,w79_115,w79_116,w79_117,w79_118,w79_119,w79_120,w79_121,w79_122,w79_123,w79_124,w79_125,w79_126,
	w80_0,w80_1,w80_2,w80_3,w80_4,w80_5,w80_6,w80_7,w80_8,w80_9,w80_10,w80_11,w80_12,w80_13,w80_14,w80_15,w80_16,
		w80_17,w80_18,w80_19,w80_20,w80_21,w80_22,w80_23,w80_24,w80_25,w80_26,w80_27,w80_28,w80_29,w80_30,w80_31,w80_32,
		w80_33,w80_34,w80_35,w80_36,w80_37,w80_38,w80_39,w80_40,w80_41,w80_42,w80_43,w80_44,w80_45,w80_46,w80_47,w80_48,
		w80_49,w80_50,w80_51,w80_52,w80_53,w80_54,w80_55,w80_56,w80_57,w80_58,w80_59,w80_60,w80_61,w80_62,w80_63,w80_64,
		w80_65,w80_66,w80_67,w80_68,w80_69,w80_70,w80_71,w80_72,w80_73,w80_74,w80_75,w80_76,w80_77,w80_78,w80_79,w80_80,
		w80_81,w80_82,w80_83,w80_84,w80_85,w80_86,w80_87,w80_88,w80_89,w80_90,w80_91,w80_92,w80_93,w80_94,w80_95,w80_96,
		w80_97,w80_98,w80_99,w80_100,w80_101,w80_102,w80_103,w80_104,w80_105,w80_106,w80_107,w80_108,w80_109,w80_110,w80_111,w80_112,
		w80_113,w80_114,w80_115,w80_116,w80_117,w80_118,w80_119,w80_120,w80_121,w80_122,w80_123,w80_124,w80_125,w80_126,
	w81_0,w81_1,w81_2,w81_3,w81_4,w81_5,w81_6,w81_7,w81_8,w81_9,w81_10,w81_11,w81_12,w81_13,w81_14,w81_15,w81_16,
		w81_17,w81_18,w81_19,w81_20,w81_21,w81_22,w81_23,w81_24,w81_25,w81_26,w81_27,w81_28,w81_29,w81_30,w81_31,w81_32,
		w81_33,w81_34,w81_35,w81_36,w81_37,w81_38,w81_39,w81_40,w81_41,w81_42,w81_43,w81_44,w81_45,w81_46,w81_47,w81_48,
		w81_49,w81_50,w81_51,w81_52,w81_53,w81_54,w81_55,w81_56,w81_57,w81_58,w81_59,w81_60,w81_61,w81_62,w81_63,w81_64,
		w81_65,w81_66,w81_67,w81_68,w81_69,w81_70,w81_71,w81_72,w81_73,w81_74,w81_75,w81_76,w81_77,w81_78,w81_79,w81_80,
		w81_81,w81_82,w81_83,w81_84,w81_85,w81_86,w81_87,w81_88,w81_89,w81_90,w81_91,w81_92,w81_93,w81_94,w81_95,w81_96,
		w81_97,w81_98,w81_99,w81_100,w81_101,w81_102,w81_103,w81_104,w81_105,w81_106,w81_107,w81_108,w81_109,w81_110,w81_111,w81_112,
		w81_113,w81_114,w81_115,w81_116,w81_117,w81_118,w81_119,w81_120,w81_121,w81_122,w81_123,w81_124,w81_125,w81_126,
	w82_0,w82_1,w82_2,w82_3,w82_4,w82_5,w82_6,w82_7,w82_8,w82_9,w82_10,w82_11,w82_12,w82_13,w82_14,w82_15,w82_16,
		w82_17,w82_18,w82_19,w82_20,w82_21,w82_22,w82_23,w82_24,w82_25,w82_26,w82_27,w82_28,w82_29,w82_30,w82_31,w82_32,
		w82_33,w82_34,w82_35,w82_36,w82_37,w82_38,w82_39,w82_40,w82_41,w82_42,w82_43,w82_44,w82_45,w82_46,w82_47,w82_48,
		w82_49,w82_50,w82_51,w82_52,w82_53,w82_54,w82_55,w82_56,w82_57,w82_58,w82_59,w82_60,w82_61,w82_62,w82_63,w82_64,
		w82_65,w82_66,w82_67,w82_68,w82_69,w82_70,w82_71,w82_72,w82_73,w82_74,w82_75,w82_76,w82_77,w82_78,w82_79,w82_80,
		w82_81,w82_82,w82_83,w82_84,w82_85,w82_86,w82_87,w82_88,w82_89,w82_90,w82_91,w82_92,w82_93,w82_94,w82_95,w82_96,
		w82_97,w82_98,w82_99,w82_100,w82_101,w82_102,w82_103,w82_104,w82_105,w82_106,w82_107,w82_108,w82_109,w82_110,w82_111,w82_112,
		w82_113,w82_114,w82_115,w82_116,w82_117,w82_118,w82_119,w82_120,w82_121,w82_122,w82_123,w82_124,w82_125,w82_126,
	w83_0,w83_1,w83_2,w83_3,w83_4,w83_5,w83_6,w83_7,w83_8,w83_9,w83_10,w83_11,w83_12,w83_13,w83_14,w83_15,w83_16,
		w83_17,w83_18,w83_19,w83_20,w83_21,w83_22,w83_23,w83_24,w83_25,w83_26,w83_27,w83_28,w83_29,w83_30,w83_31,w83_32,
		w83_33,w83_34,w83_35,w83_36,w83_37,w83_38,w83_39,w83_40,w83_41,w83_42,w83_43,w83_44,w83_45,w83_46,w83_47,w83_48,
		w83_49,w83_50,w83_51,w83_52,w83_53,w83_54,w83_55,w83_56,w83_57,w83_58,w83_59,w83_60,w83_61,w83_62,w83_63,w83_64,
		w83_65,w83_66,w83_67,w83_68,w83_69,w83_70,w83_71,w83_72,w83_73,w83_74,w83_75,w83_76,w83_77,w83_78,w83_79,w83_80,
		w83_81,w83_82,w83_83,w83_84,w83_85,w83_86,w83_87,w83_88,w83_89,w83_90,w83_91,w83_92,w83_93,w83_94,w83_95,w83_96,
		w83_97,w83_98,w83_99,w83_100,w83_101,w83_102,w83_103,w83_104,w83_105,w83_106,w83_107,w83_108,w83_109,w83_110,w83_111,w83_112,
		w83_113,w83_114,w83_115,w83_116,w83_117,w83_118,w83_119,w83_120,w83_121,w83_122,w83_123,w83_124,w83_125,w83_126,
	w84_0,w84_1,w84_2,w84_3,w84_4,w84_5,w84_6,w84_7,w84_8,w84_9,w84_10,w84_11,w84_12,w84_13,w84_14,w84_15,w84_16,
		w84_17,w84_18,w84_19,w84_20,w84_21,w84_22,w84_23,w84_24,w84_25,w84_26,w84_27,w84_28,w84_29,w84_30,w84_31,w84_32,
		w84_33,w84_34,w84_35,w84_36,w84_37,w84_38,w84_39,w84_40,w84_41,w84_42,w84_43,w84_44,w84_45,w84_46,w84_47,w84_48,
		w84_49,w84_50,w84_51,w84_52,w84_53,w84_54,w84_55,w84_56,w84_57,w84_58,w84_59,w84_60,w84_61,w84_62,w84_63,w84_64,
		w84_65,w84_66,w84_67,w84_68,w84_69,w84_70,w84_71,w84_72,w84_73,w84_74,w84_75,w84_76,w84_77,w84_78,w84_79,w84_80,
		w84_81,w84_82,w84_83,w84_84,w84_85,w84_86,w84_87,w84_88,w84_89,w84_90,w84_91,w84_92,w84_93,w84_94,w84_95,w84_96,
		w84_97,w84_98,w84_99,w84_100,w84_101,w84_102,w84_103,w84_104,w84_105,w84_106,w84_107,w84_108,w84_109,w84_110,w84_111,w84_112,
		w84_113,w84_114,w84_115,w84_116,w84_117,w84_118,w84_119,w84_120,w84_121,w84_122,w84_123,w84_124,w84_125,w84_126,
	w85_0,w85_1,w85_2,w85_3,w85_4,w85_5,w85_6,w85_7,w85_8,w85_9,w85_10,w85_11,w85_12,w85_13,w85_14,w85_15,w85_16,
		w85_17,w85_18,w85_19,w85_20,w85_21,w85_22,w85_23,w85_24,w85_25,w85_26,w85_27,w85_28,w85_29,w85_30,w85_31,w85_32,
		w85_33,w85_34,w85_35,w85_36,w85_37,w85_38,w85_39,w85_40,w85_41,w85_42,w85_43,w85_44,w85_45,w85_46,w85_47,w85_48,
		w85_49,w85_50,w85_51,w85_52,w85_53,w85_54,w85_55,w85_56,w85_57,w85_58,w85_59,w85_60,w85_61,w85_62,w85_63,w85_64,
		w85_65,w85_66,w85_67,w85_68,w85_69,w85_70,w85_71,w85_72,w85_73,w85_74,w85_75,w85_76,w85_77,w85_78,w85_79,w85_80,
		w85_81,w85_82,w85_83,w85_84,w85_85,w85_86,w85_87,w85_88,w85_89,w85_90,w85_91,w85_92,w85_93,w85_94,w85_95,w85_96,
		w85_97,w85_98,w85_99,w85_100,w85_101,w85_102,w85_103,w85_104,w85_105,w85_106,w85_107,w85_108,w85_109,w85_110,w85_111,w85_112,
		w85_113,w85_114,w85_115,w85_116,w85_117,w85_118,w85_119,w85_120,w85_121,w85_122,w85_123,w85_124,w85_125,w85_126,
	w86_0,w86_1,w86_2,w86_3,w86_4,w86_5,w86_6,w86_7,w86_8,w86_9,w86_10,w86_11,w86_12,w86_13,w86_14,w86_15,w86_16,
		w86_17,w86_18,w86_19,w86_20,w86_21,w86_22,w86_23,w86_24,w86_25,w86_26,w86_27,w86_28,w86_29,w86_30,w86_31,w86_32,
		w86_33,w86_34,w86_35,w86_36,w86_37,w86_38,w86_39,w86_40,w86_41,w86_42,w86_43,w86_44,w86_45,w86_46,w86_47,w86_48,
		w86_49,w86_50,w86_51,w86_52,w86_53,w86_54,w86_55,w86_56,w86_57,w86_58,w86_59,w86_60,w86_61,w86_62,w86_63,w86_64,
		w86_65,w86_66,w86_67,w86_68,w86_69,w86_70,w86_71,w86_72,w86_73,w86_74,w86_75,w86_76,w86_77,w86_78,w86_79,w86_80,
		w86_81,w86_82,w86_83,w86_84,w86_85,w86_86,w86_87,w86_88,w86_89,w86_90,w86_91,w86_92,w86_93,w86_94,w86_95,w86_96,
		w86_97,w86_98,w86_99,w86_100,w86_101,w86_102,w86_103,w86_104,w86_105,w86_106,w86_107,w86_108,w86_109,w86_110,w86_111,w86_112,
		w86_113,w86_114,w86_115,w86_116,w86_117,w86_118,w86_119,w86_120,w86_121,w86_122,w86_123,w86_124,w86_125,w86_126,
	w87_0,w87_1,w87_2,w87_3,w87_4,w87_5,w87_6,w87_7,w87_8,w87_9,w87_10,w87_11,w87_12,w87_13,w87_14,w87_15,w87_16,
		w87_17,w87_18,w87_19,w87_20,w87_21,w87_22,w87_23,w87_24,w87_25,w87_26,w87_27,w87_28,w87_29,w87_30,w87_31,w87_32,
		w87_33,w87_34,w87_35,w87_36,w87_37,w87_38,w87_39,w87_40,w87_41,w87_42,w87_43,w87_44,w87_45,w87_46,w87_47,w87_48,
		w87_49,w87_50,w87_51,w87_52,w87_53,w87_54,w87_55,w87_56,w87_57,w87_58,w87_59,w87_60,w87_61,w87_62,w87_63,w87_64,
		w87_65,w87_66,w87_67,w87_68,w87_69,w87_70,w87_71,w87_72,w87_73,w87_74,w87_75,w87_76,w87_77,w87_78,w87_79,w87_80,
		w87_81,w87_82,w87_83,w87_84,w87_85,w87_86,w87_87,w87_88,w87_89,w87_90,w87_91,w87_92,w87_93,w87_94,w87_95,w87_96,
		w87_97,w87_98,w87_99,w87_100,w87_101,w87_102,w87_103,w87_104,w87_105,w87_106,w87_107,w87_108,w87_109,w87_110,w87_111,w87_112,
		w87_113,w87_114,w87_115,w87_116,w87_117,w87_118,w87_119,w87_120,w87_121,w87_122,w87_123,w87_124,w87_125,w87_126,
	w88_0,w88_1,w88_2,w88_3,w88_4,w88_5,w88_6,w88_7,w88_8,w88_9,w88_10,w88_11,w88_12,w88_13,w88_14,w88_15,w88_16,
		w88_17,w88_18,w88_19,w88_20,w88_21,w88_22,w88_23,w88_24,w88_25,w88_26,w88_27,w88_28,w88_29,w88_30,w88_31,w88_32,
		w88_33,w88_34,w88_35,w88_36,w88_37,w88_38,w88_39,w88_40,w88_41,w88_42,w88_43,w88_44,w88_45,w88_46,w88_47,w88_48,
		w88_49,w88_50,w88_51,w88_52,w88_53,w88_54,w88_55,w88_56,w88_57,w88_58,w88_59,w88_60,w88_61,w88_62,w88_63,w88_64,
		w88_65,w88_66,w88_67,w88_68,w88_69,w88_70,w88_71,w88_72,w88_73,w88_74,w88_75,w88_76,w88_77,w88_78,w88_79,w88_80,
		w88_81,w88_82,w88_83,w88_84,w88_85,w88_86,w88_87,w88_88,w88_89,w88_90,w88_91,w88_92,w88_93,w88_94,w88_95,w88_96,
		w88_97,w88_98,w88_99,w88_100,w88_101,w88_102,w88_103,w88_104,w88_105,w88_106,w88_107,w88_108,w88_109,w88_110,w88_111,w88_112,
		w88_113,w88_114,w88_115,w88_116,w88_117,w88_118,w88_119,w88_120,w88_121,w88_122,w88_123,w88_124,w88_125,w88_126,
	w89_0,w89_1,w89_2,w89_3,w89_4,w89_5,w89_6,w89_7,w89_8,w89_9,w89_10,w89_11,w89_12,w89_13,w89_14,w89_15,w89_16,
		w89_17,w89_18,w89_19,w89_20,w89_21,w89_22,w89_23,w89_24,w89_25,w89_26,w89_27,w89_28,w89_29,w89_30,w89_31,w89_32,
		w89_33,w89_34,w89_35,w89_36,w89_37,w89_38,w89_39,w89_40,w89_41,w89_42,w89_43,w89_44,w89_45,w89_46,w89_47,w89_48,
		w89_49,w89_50,w89_51,w89_52,w89_53,w89_54,w89_55,w89_56,w89_57,w89_58,w89_59,w89_60,w89_61,w89_62,w89_63,w89_64,
		w89_65,w89_66,w89_67,w89_68,w89_69,w89_70,w89_71,w89_72,w89_73,w89_74,w89_75,w89_76,w89_77,w89_78,w89_79,w89_80,
		w89_81,w89_82,w89_83,w89_84,w89_85,w89_86,w89_87,w89_88,w89_89,w89_90,w89_91,w89_92,w89_93,w89_94,w89_95,w89_96,
		w89_97,w89_98,w89_99,w89_100,w89_101,w89_102,w89_103,w89_104,w89_105,w89_106,w89_107,w89_108,w89_109,w89_110,w89_111,w89_112,
		w89_113,w89_114,w89_115,w89_116,w89_117,w89_118,w89_119,w89_120,w89_121,w89_122,w89_123,w89_124,w89_125,w89_126,
	w90_0,w90_1,w90_2,w90_3,w90_4,w90_5,w90_6,w90_7,w90_8,w90_9,w90_10,w90_11,w90_12,w90_13,w90_14,w90_15,w90_16,
		w90_17,w90_18,w90_19,w90_20,w90_21,w90_22,w90_23,w90_24,w90_25,w90_26,w90_27,w90_28,w90_29,w90_30,w90_31,w90_32,
		w90_33,w90_34,w90_35,w90_36,w90_37,w90_38,w90_39,w90_40,w90_41,w90_42,w90_43,w90_44,w90_45,w90_46,w90_47,w90_48,
		w90_49,w90_50,w90_51,w90_52,w90_53,w90_54,w90_55,w90_56,w90_57,w90_58,w90_59,w90_60,w90_61,w90_62,w90_63,w90_64,
		w90_65,w90_66,w90_67,w90_68,w90_69,w90_70,w90_71,w90_72,w90_73,w90_74,w90_75,w90_76,w90_77,w90_78,w90_79,w90_80,
		w90_81,w90_82,w90_83,w90_84,w90_85,w90_86,w90_87,w90_88,w90_89,w90_90,w90_91,w90_92,w90_93,w90_94,w90_95,w90_96,
		w90_97,w90_98,w90_99,w90_100,w90_101,w90_102,w90_103,w90_104,w90_105,w90_106,w90_107,w90_108,w90_109,w90_110,w90_111,w90_112,
		w90_113,w90_114,w90_115,w90_116,w90_117,w90_118,w90_119,w90_120,w90_121,w90_122,w90_123,w90_124,w90_125,w90_126,
	w91_0,w91_1,w91_2,w91_3,w91_4,w91_5,w91_6,w91_7,w91_8,w91_9,w91_10,w91_11,w91_12,w91_13,w91_14,w91_15,w91_16,
		w91_17,w91_18,w91_19,w91_20,w91_21,w91_22,w91_23,w91_24,w91_25,w91_26,w91_27,w91_28,w91_29,w91_30,w91_31,w91_32,
		w91_33,w91_34,w91_35,w91_36,w91_37,w91_38,w91_39,w91_40,w91_41,w91_42,w91_43,w91_44,w91_45,w91_46,w91_47,w91_48,
		w91_49,w91_50,w91_51,w91_52,w91_53,w91_54,w91_55,w91_56,w91_57,w91_58,w91_59,w91_60,w91_61,w91_62,w91_63,w91_64,
		w91_65,w91_66,w91_67,w91_68,w91_69,w91_70,w91_71,w91_72,w91_73,w91_74,w91_75,w91_76,w91_77,w91_78,w91_79,w91_80,
		w91_81,w91_82,w91_83,w91_84,w91_85,w91_86,w91_87,w91_88,w91_89,w91_90,w91_91,w91_92,w91_93,w91_94,w91_95,w91_96,
		w91_97,w91_98,w91_99,w91_100,w91_101,w91_102,w91_103,w91_104,w91_105,w91_106,w91_107,w91_108,w91_109,w91_110,w91_111,w91_112,
		w91_113,w91_114,w91_115,w91_116,w91_117,w91_118,w91_119,w91_120,w91_121,w91_122,w91_123,w91_124,w91_125,w91_126,
	w92_0,w92_1,w92_2,w92_3,w92_4,w92_5,w92_6,w92_7,w92_8,w92_9,w92_10,w92_11,w92_12,w92_13,w92_14,w92_15,w92_16,
		w92_17,w92_18,w92_19,w92_20,w92_21,w92_22,w92_23,w92_24,w92_25,w92_26,w92_27,w92_28,w92_29,w92_30,w92_31,w92_32,
		w92_33,w92_34,w92_35,w92_36,w92_37,w92_38,w92_39,w92_40,w92_41,w92_42,w92_43,w92_44,w92_45,w92_46,w92_47,w92_48,
		w92_49,w92_50,w92_51,w92_52,w92_53,w92_54,w92_55,w92_56,w92_57,w92_58,w92_59,w92_60,w92_61,w92_62,w92_63,w92_64,
		w92_65,w92_66,w92_67,w92_68,w92_69,w92_70,w92_71,w92_72,w92_73,w92_74,w92_75,w92_76,w92_77,w92_78,w92_79,w92_80,
		w92_81,w92_82,w92_83,w92_84,w92_85,w92_86,w92_87,w92_88,w92_89,w92_90,w92_91,w92_92,w92_93,w92_94,w92_95,w92_96,
		w92_97,w92_98,w92_99,w92_100,w92_101,w92_102,w92_103,w92_104,w92_105,w92_106,w92_107,w92_108,w92_109,w92_110,w92_111,w92_112,
		w92_113,w92_114,w92_115,w92_116,w92_117,w92_118,w92_119,w92_120,w92_121,w92_122,w92_123,w92_124,w92_125,w92_126,
	w93_0,w93_1,w93_2,w93_3,w93_4,w93_5,w93_6,w93_7,w93_8,w93_9,w93_10,w93_11,w93_12,w93_13,w93_14,w93_15,w93_16,
		w93_17,w93_18,w93_19,w93_20,w93_21,w93_22,w93_23,w93_24,w93_25,w93_26,w93_27,w93_28,w93_29,w93_30,w93_31,w93_32,
		w93_33,w93_34,w93_35,w93_36,w93_37,w93_38,w93_39,w93_40,w93_41,w93_42,w93_43,w93_44,w93_45,w93_46,w93_47,w93_48,
		w93_49,w93_50,w93_51,w93_52,w93_53,w93_54,w93_55,w93_56,w93_57,w93_58,w93_59,w93_60,w93_61,w93_62,w93_63,w93_64,
		w93_65,w93_66,w93_67,w93_68,w93_69,w93_70,w93_71,w93_72,w93_73,w93_74,w93_75,w93_76,w93_77,w93_78,w93_79,w93_80,
		w93_81,w93_82,w93_83,w93_84,w93_85,w93_86,w93_87,w93_88,w93_89,w93_90,w93_91,w93_92,w93_93,w93_94,w93_95,w93_96,
		w93_97,w93_98,w93_99,w93_100,w93_101,w93_102,w93_103,w93_104,w93_105,w93_106,w93_107,w93_108,w93_109,w93_110,w93_111,w93_112,
		w93_113,w93_114,w93_115,w93_116,w93_117,w93_118,w93_119,w93_120,w93_121,w93_122,w93_123,w93_124,w93_125,w93_126,
	w94_0,w94_1,w94_2,w94_3,w94_4,w94_5,w94_6,w94_7,w94_8,w94_9,w94_10,w94_11,w94_12,w94_13,w94_14,w94_15,w94_16,
		w94_17,w94_18,w94_19,w94_20,w94_21,w94_22,w94_23,w94_24,w94_25,w94_26,w94_27,w94_28,w94_29,w94_30,w94_31,w94_32,
		w94_33,w94_34,w94_35,w94_36,w94_37,w94_38,w94_39,w94_40,w94_41,w94_42,w94_43,w94_44,w94_45,w94_46,w94_47,w94_48,
		w94_49,w94_50,w94_51,w94_52,w94_53,w94_54,w94_55,w94_56,w94_57,w94_58,w94_59,w94_60,w94_61,w94_62,w94_63,w94_64,
		w94_65,w94_66,w94_67,w94_68,w94_69,w94_70,w94_71,w94_72,w94_73,w94_74,w94_75,w94_76,w94_77,w94_78,w94_79,w94_80,
		w94_81,w94_82,w94_83,w94_84,w94_85,w94_86,w94_87,w94_88,w94_89,w94_90,w94_91,w94_92,w94_93,w94_94,w94_95,w94_96,
		w94_97,w94_98,w94_99,w94_100,w94_101,w94_102,w94_103,w94_104,w94_105,w94_106,w94_107,w94_108,w94_109,w94_110,w94_111,w94_112,
		w94_113,w94_114,w94_115,w94_116,w94_117,w94_118,w94_119,w94_120,w94_121,w94_122,w94_123,w94_124,w94_125,w94_126,
	w95_0,w95_1,w95_2,w95_3,w95_4,w95_5,w95_6,w95_7,w95_8,w95_9,w95_10,w95_11,w95_12,w95_13,w95_14,w95_15,w95_16,
		w95_17,w95_18,w95_19,w95_20,w95_21,w95_22,w95_23,w95_24,w95_25,w95_26,w95_27,w95_28,w95_29,w95_30,w95_31,w95_32,
		w95_33,w95_34,w95_35,w95_36,w95_37,w95_38,w95_39,w95_40,w95_41,w95_42,w95_43,w95_44,w95_45,w95_46,w95_47,w95_48,
		w95_49,w95_50,w95_51,w95_52,w95_53,w95_54,w95_55,w95_56,w95_57,w95_58,w95_59,w95_60,w95_61,w95_62,w95_63,w95_64,
		w95_65,w95_66,w95_67,w95_68,w95_69,w95_70,w95_71,w95_72,w95_73,w95_74,w95_75,w95_76,w95_77,w95_78,w95_79,w95_80,
		w95_81,w95_82,w95_83,w95_84,w95_85,w95_86,w95_87,w95_88,w95_89,w95_90,w95_91,w95_92,w95_93,w95_94,w95_95,w95_96,
		w95_97,w95_98,w95_99,w95_100,w95_101,w95_102,w95_103,w95_104,w95_105,w95_106,w95_107,w95_108,w95_109,w95_110,w95_111,w95_112,
		w95_113,w95_114,w95_115,w95_116,w95_117,w95_118,w95_119,w95_120,w95_121,w95_122,w95_123,w95_124,w95_125,w95_126,
	w96_0,w96_1,w96_2,w96_3,w96_4,w96_5,w96_6,w96_7,w96_8,w96_9,w96_10,w96_11,w96_12,w96_13,w96_14,w96_15,w96_16,
		w96_17,w96_18,w96_19,w96_20,w96_21,w96_22,w96_23,w96_24,w96_25,w96_26,w96_27,w96_28,w96_29,w96_30,w96_31,w96_32,
		w96_33,w96_34,w96_35,w96_36,w96_37,w96_38,w96_39,w96_40,w96_41,w96_42,w96_43,w96_44,w96_45,w96_46,w96_47,w96_48,
		w96_49,w96_50,w96_51,w96_52,w96_53,w96_54,w96_55,w96_56,w96_57,w96_58,w96_59,w96_60,w96_61,w96_62,w96_63,w96_64,
		w96_65,w96_66,w96_67,w96_68,w96_69,w96_70,w96_71,w96_72,w96_73,w96_74,w96_75,w96_76,w96_77,w96_78,w96_79,w96_80,
		w96_81,w96_82,w96_83,w96_84,w96_85,w96_86,w96_87,w96_88,w96_89,w96_90,w96_91,w96_92,w96_93,w96_94,w96_95,w96_96,
		w96_97,w96_98,w96_99,w96_100,w96_101,w96_102,w96_103,w96_104,w96_105,w96_106,w96_107,w96_108,w96_109,w96_110,w96_111,w96_112,
		w96_113,w96_114,w96_115,w96_116,w96_117,w96_118,w96_119,w96_120,w96_121,w96_122,w96_123,w96_124,w96_125,w96_126,
	w97_0,w97_1,w97_2,w97_3,w97_4,w97_5,w97_6,w97_7,w97_8,w97_9,w97_10,w97_11,w97_12,w97_13,w97_14,w97_15,w97_16,
		w97_17,w97_18,w97_19,w97_20,w97_21,w97_22,w97_23,w97_24,w97_25,w97_26,w97_27,w97_28,w97_29,w97_30,w97_31,w97_32,
		w97_33,w97_34,w97_35,w97_36,w97_37,w97_38,w97_39,w97_40,w97_41,w97_42,w97_43,w97_44,w97_45,w97_46,w97_47,w97_48,
		w97_49,w97_50,w97_51,w97_52,w97_53,w97_54,w97_55,w97_56,w97_57,w97_58,w97_59,w97_60,w97_61,w97_62,w97_63,w97_64,
		w97_65,w97_66,w97_67,w97_68,w97_69,w97_70,w97_71,w97_72,w97_73,w97_74,w97_75,w97_76,w97_77,w97_78,w97_79,w97_80,
		w97_81,w97_82,w97_83,w97_84,w97_85,w97_86,w97_87,w97_88,w97_89,w97_90,w97_91,w97_92,w97_93,w97_94,w97_95,w97_96,
		w97_97,w97_98,w97_99,w97_100,w97_101,w97_102,w97_103,w97_104,w97_105,w97_106,w97_107,w97_108,w97_109,w97_110,w97_111,w97_112,
		w97_113,w97_114,w97_115,w97_116,w97_117,w97_118,w97_119,w97_120,w97_121,w97_122,w97_123,w97_124,w97_125,w97_126,
	w98_0,w98_1,w98_2,w98_3,w98_4,w98_5,w98_6,w98_7,w98_8,w98_9,w98_10,w98_11,w98_12,w98_13,w98_14,w98_15,w98_16,
		w98_17,w98_18,w98_19,w98_20,w98_21,w98_22,w98_23,w98_24,w98_25,w98_26,w98_27,w98_28,w98_29,w98_30,w98_31,w98_32,
		w98_33,w98_34,w98_35,w98_36,w98_37,w98_38,w98_39,w98_40,w98_41,w98_42,w98_43,w98_44,w98_45,w98_46,w98_47,w98_48,
		w98_49,w98_50,w98_51,w98_52,w98_53,w98_54,w98_55,w98_56,w98_57,w98_58,w98_59,w98_60,w98_61,w98_62,w98_63,w98_64,
		w98_65,w98_66,w98_67,w98_68,w98_69,w98_70,w98_71,w98_72,w98_73,w98_74,w98_75,w98_76,w98_77,w98_78,w98_79,w98_80,
		w98_81,w98_82,w98_83,w98_84,w98_85,w98_86,w98_87,w98_88,w98_89,w98_90,w98_91,w98_92,w98_93,w98_94,w98_95,w98_96,
		w98_97,w98_98,w98_99,w98_100,w98_101,w98_102,w98_103,w98_104,w98_105,w98_106,w98_107,w98_108,w98_109,w98_110,w98_111,w98_112,
		w98_113,w98_114,w98_115,w98_116,w98_117,w98_118,w98_119,w98_120,w98_121,w98_122,w98_123,w98_124,w98_125,w98_126,
	w99_0,w99_1,w99_2,w99_3,w99_4,w99_5,w99_6,w99_7,w99_8,w99_9,w99_10,w99_11,w99_12,w99_13,w99_14,w99_15,w99_16,
		w99_17,w99_18,w99_19,w99_20,w99_21,w99_22,w99_23,w99_24,w99_25,w99_26,w99_27,w99_28,w99_29,w99_30,w99_31,w99_32,
		w99_33,w99_34,w99_35,w99_36,w99_37,w99_38,w99_39,w99_40,w99_41,w99_42,w99_43,w99_44,w99_45,w99_46,w99_47,w99_48,
		w99_49,w99_50,w99_51,w99_52,w99_53,w99_54,w99_55,w99_56,w99_57,w99_58,w99_59,w99_60,w99_61,w99_62,w99_63,w99_64,
		w99_65,w99_66,w99_67,w99_68,w99_69,w99_70,w99_71,w99_72,w99_73,w99_74,w99_75,w99_76,w99_77,w99_78,w99_79,w99_80,
		w99_81,w99_82,w99_83,w99_84,w99_85,w99_86,w99_87,w99_88,w99_89,w99_90,w99_91,w99_92,w99_93,w99_94,w99_95,w99_96,
		w99_97,w99_98,w99_99,w99_100,w99_101,w99_102,w99_103,w99_104,w99_105,w99_106,w99_107,w99_108,w99_109,w99_110,w99_111,w99_112,
		w99_113,w99_114,w99_115,w99_116,w99_117,w99_118,w99_119,w99_120,w99_121,w99_122,w99_123,w99_124,w99_125,w99_126,
	w100_0,w100_1,w100_2,w100_3,w100_4,w100_5,w100_6,w100_7,w100_8,w100_9,w100_10,w100_11,w100_12,w100_13,w100_14,w100_15,w100_16,
		w100_17,w100_18,w100_19,w100_20,w100_21,w100_22,w100_23,w100_24,w100_25,w100_26,w100_27,w100_28,w100_29,w100_30,w100_31,w100_32,
		w100_33,w100_34,w100_35,w100_36,w100_37,w100_38,w100_39,w100_40,w100_41,w100_42,w100_43,w100_44,w100_45,w100_46,w100_47,w100_48,
		w100_49,w100_50,w100_51,w100_52,w100_53,w100_54,w100_55,w100_56,w100_57,w100_58,w100_59,w100_60,w100_61,w100_62,w100_63,w100_64,
		w100_65,w100_66,w100_67,w100_68,w100_69,w100_70,w100_71,w100_72,w100_73,w100_74,w100_75,w100_76,w100_77,w100_78,w100_79,w100_80,
		w100_81,w100_82,w100_83,w100_84,w100_85,w100_86,w100_87,w100_88,w100_89,w100_90,w100_91,w100_92,w100_93,w100_94,w100_95,w100_96,
		w100_97,w100_98,w100_99,w100_100,w100_101,w100_102,w100_103,w100_104,w100_105,w100_106,w100_107,w100_108,w100_109,w100_110,w100_111,w100_112,
		w100_113,w100_114,w100_115,w100_116,w100_117,w100_118,w100_119,w100_120,w100_121,w100_122,w100_123,w100_124,w100_125,w100_126,
	w101_0,w101_1,w101_2,w101_3,w101_4,w101_5,w101_6,w101_7,w101_8,w101_9,w101_10,w101_11,w101_12,w101_13,w101_14,w101_15,w101_16,
		w101_17,w101_18,w101_19,w101_20,w101_21,w101_22,w101_23,w101_24,w101_25,w101_26,w101_27,w101_28,w101_29,w101_30,w101_31,w101_32,
		w101_33,w101_34,w101_35,w101_36,w101_37,w101_38,w101_39,w101_40,w101_41,w101_42,w101_43,w101_44,w101_45,w101_46,w101_47,w101_48,
		w101_49,w101_50,w101_51,w101_52,w101_53,w101_54,w101_55,w101_56,w101_57,w101_58,w101_59,w101_60,w101_61,w101_62,w101_63,w101_64,
		w101_65,w101_66,w101_67,w101_68,w101_69,w101_70,w101_71,w101_72,w101_73,w101_74,w101_75,w101_76,w101_77,w101_78,w101_79,w101_80,
		w101_81,w101_82,w101_83,w101_84,w101_85,w101_86,w101_87,w101_88,w101_89,w101_90,w101_91,w101_92,w101_93,w101_94,w101_95,w101_96,
		w101_97,w101_98,w101_99,w101_100,w101_101,w101_102,w101_103,w101_104,w101_105,w101_106,w101_107,w101_108,w101_109,w101_110,w101_111,w101_112,
		w101_113,w101_114,w101_115,w101_116,w101_117,w101_118,w101_119,w101_120,w101_121,w101_122,w101_123,w101_124,w101_125,w101_126,
	w102_0,w102_1,w102_2,w102_3,w102_4,w102_5,w102_6,w102_7,w102_8,w102_9,w102_10,w102_11,w102_12,w102_13,w102_14,w102_15,w102_16,
		w102_17,w102_18,w102_19,w102_20,w102_21,w102_22,w102_23,w102_24,w102_25,w102_26,w102_27,w102_28,w102_29,w102_30,w102_31,w102_32,
		w102_33,w102_34,w102_35,w102_36,w102_37,w102_38,w102_39,w102_40,w102_41,w102_42,w102_43,w102_44,w102_45,w102_46,w102_47,w102_48,
		w102_49,w102_50,w102_51,w102_52,w102_53,w102_54,w102_55,w102_56,w102_57,w102_58,w102_59,w102_60,w102_61,w102_62,w102_63,w102_64,
		w102_65,w102_66,w102_67,w102_68,w102_69,w102_70,w102_71,w102_72,w102_73,w102_74,w102_75,w102_76,w102_77,w102_78,w102_79,w102_80,
		w102_81,w102_82,w102_83,w102_84,w102_85,w102_86,w102_87,w102_88,w102_89,w102_90,w102_91,w102_92,w102_93,w102_94,w102_95,w102_96,
		w102_97,w102_98,w102_99,w102_100,w102_101,w102_102,w102_103,w102_104,w102_105,w102_106,w102_107,w102_108,w102_109,w102_110,w102_111,w102_112,
		w102_113,w102_114,w102_115,w102_116,w102_117,w102_118,w102_119,w102_120,w102_121,w102_122,w102_123,w102_124,w102_125,w102_126,
	w103_0,w103_1,w103_2,w103_3,w103_4,w103_5,w103_6,w103_7,w103_8,w103_9,w103_10,w103_11,w103_12,w103_13,w103_14,w103_15,w103_16,
		w103_17,w103_18,w103_19,w103_20,w103_21,w103_22,w103_23,w103_24,w103_25,w103_26,w103_27,w103_28,w103_29,w103_30,w103_31,w103_32,
		w103_33,w103_34,w103_35,w103_36,w103_37,w103_38,w103_39,w103_40,w103_41,w103_42,w103_43,w103_44,w103_45,w103_46,w103_47,w103_48,
		w103_49,w103_50,w103_51,w103_52,w103_53,w103_54,w103_55,w103_56,w103_57,w103_58,w103_59,w103_60,w103_61,w103_62,w103_63,w103_64,
		w103_65,w103_66,w103_67,w103_68,w103_69,w103_70,w103_71,w103_72,w103_73,w103_74,w103_75,w103_76,w103_77,w103_78,w103_79,w103_80,
		w103_81,w103_82,w103_83,w103_84,w103_85,w103_86,w103_87,w103_88,w103_89,w103_90,w103_91,w103_92,w103_93,w103_94,w103_95,w103_96,
		w103_97,w103_98,w103_99,w103_100,w103_101,w103_102,w103_103,w103_104,w103_105,w103_106,w103_107,w103_108,w103_109,w103_110,w103_111,w103_112,
		w103_113,w103_114,w103_115,w103_116,w103_117,w103_118,w103_119,w103_120,w103_121,w103_122,w103_123,w103_124,w103_125,w103_126,
	w104_0,w104_1,w104_2,w104_3,w104_4,w104_5,w104_6,w104_7,w104_8,w104_9,w104_10,w104_11,w104_12,w104_13,w104_14,w104_15,w104_16,
		w104_17,w104_18,w104_19,w104_20,w104_21,w104_22,w104_23,w104_24,w104_25,w104_26,w104_27,w104_28,w104_29,w104_30,w104_31,w104_32,
		w104_33,w104_34,w104_35,w104_36,w104_37,w104_38,w104_39,w104_40,w104_41,w104_42,w104_43,w104_44,w104_45,w104_46,w104_47,w104_48,
		w104_49,w104_50,w104_51,w104_52,w104_53,w104_54,w104_55,w104_56,w104_57,w104_58,w104_59,w104_60,w104_61,w104_62,w104_63,w104_64,
		w104_65,w104_66,w104_67,w104_68,w104_69,w104_70,w104_71,w104_72,w104_73,w104_74,w104_75,w104_76,w104_77,w104_78,w104_79,w104_80,
		w104_81,w104_82,w104_83,w104_84,w104_85,w104_86,w104_87,w104_88,w104_89,w104_90,w104_91,w104_92,w104_93,w104_94,w104_95,w104_96,
		w104_97,w104_98,w104_99,w104_100,w104_101,w104_102,w104_103,w104_104,w104_105,w104_106,w104_107,w104_108,w104_109,w104_110,w104_111,w104_112,
		w104_113,w104_114,w104_115,w104_116,w104_117,w104_118,w104_119,w104_120,w104_121,w104_122,w104_123,w104_124,w104_125,w104_126,
	w105_0,w105_1,w105_2,w105_3,w105_4,w105_5,w105_6,w105_7,w105_8,w105_9,w105_10,w105_11,w105_12,w105_13,w105_14,w105_15,w105_16,
		w105_17,w105_18,w105_19,w105_20,w105_21,w105_22,w105_23,w105_24,w105_25,w105_26,w105_27,w105_28,w105_29,w105_30,w105_31,w105_32,
		w105_33,w105_34,w105_35,w105_36,w105_37,w105_38,w105_39,w105_40,w105_41,w105_42,w105_43,w105_44,w105_45,w105_46,w105_47,w105_48,
		w105_49,w105_50,w105_51,w105_52,w105_53,w105_54,w105_55,w105_56,w105_57,w105_58,w105_59,w105_60,w105_61,w105_62,w105_63,w105_64,
		w105_65,w105_66,w105_67,w105_68,w105_69,w105_70,w105_71,w105_72,w105_73,w105_74,w105_75,w105_76,w105_77,w105_78,w105_79,w105_80,
		w105_81,w105_82,w105_83,w105_84,w105_85,w105_86,w105_87,w105_88,w105_89,w105_90,w105_91,w105_92,w105_93,w105_94,w105_95,w105_96,
		w105_97,w105_98,w105_99,w105_100,w105_101,w105_102,w105_103,w105_104,w105_105,w105_106,w105_107,w105_108,w105_109,w105_110,w105_111,w105_112,
		w105_113,w105_114,w105_115,w105_116,w105_117,w105_118,w105_119,w105_120,w105_121,w105_122,w105_123,w105_124,w105_125,w105_126,
	w106_0,w106_1,w106_2,w106_3,w106_4,w106_5,w106_6,w106_7,w106_8,w106_9,w106_10,w106_11,w106_12,w106_13,w106_14,w106_15,w106_16,
		w106_17,w106_18,w106_19,w106_20,w106_21,w106_22,w106_23,w106_24,w106_25,w106_26,w106_27,w106_28,w106_29,w106_30,w106_31,w106_32,
		w106_33,w106_34,w106_35,w106_36,w106_37,w106_38,w106_39,w106_40,w106_41,w106_42,w106_43,w106_44,w106_45,w106_46,w106_47,w106_48,
		w106_49,w106_50,w106_51,w106_52,w106_53,w106_54,w106_55,w106_56,w106_57,w106_58,w106_59,w106_60,w106_61,w106_62,w106_63,w106_64,
		w106_65,w106_66,w106_67,w106_68,w106_69,w106_70,w106_71,w106_72,w106_73,w106_74,w106_75,w106_76,w106_77,w106_78,w106_79,w106_80,
		w106_81,w106_82,w106_83,w106_84,w106_85,w106_86,w106_87,w106_88,w106_89,w106_90,w106_91,w106_92,w106_93,w106_94,w106_95,w106_96,
		w106_97,w106_98,w106_99,w106_100,w106_101,w106_102,w106_103,w106_104,w106_105,w106_106,w106_107,w106_108,w106_109,w106_110,w106_111,w106_112,
		w106_113,w106_114,w106_115,w106_116,w106_117,w106_118,w106_119,w106_120,w106_121,w106_122,w106_123,w106_124,w106_125,w106_126,
	w107_0,w107_1,w107_2,w107_3,w107_4,w107_5,w107_6,w107_7,w107_8,w107_9,w107_10,w107_11,w107_12,w107_13,w107_14,w107_15,w107_16,
		w107_17,w107_18,w107_19,w107_20,w107_21,w107_22,w107_23,w107_24,w107_25,w107_26,w107_27,w107_28,w107_29,w107_30,w107_31,w107_32,
		w107_33,w107_34,w107_35,w107_36,w107_37,w107_38,w107_39,w107_40,w107_41,w107_42,w107_43,w107_44,w107_45,w107_46,w107_47,w107_48,
		w107_49,w107_50,w107_51,w107_52,w107_53,w107_54,w107_55,w107_56,w107_57,w107_58,w107_59,w107_60,w107_61,w107_62,w107_63,w107_64,
		w107_65,w107_66,w107_67,w107_68,w107_69,w107_70,w107_71,w107_72,w107_73,w107_74,w107_75,w107_76,w107_77,w107_78,w107_79,w107_80,
		w107_81,w107_82,w107_83,w107_84,w107_85,w107_86,w107_87,w107_88,w107_89,w107_90,w107_91,w107_92,w107_93,w107_94,w107_95,w107_96,
		w107_97,w107_98,w107_99,w107_100,w107_101,w107_102,w107_103,w107_104,w107_105,w107_106,w107_107,w107_108,w107_109,w107_110,w107_111,w107_112,
		w107_113,w107_114,w107_115,w107_116,w107_117,w107_118,w107_119,w107_120,w107_121,w107_122,w107_123,w107_124,w107_125,w107_126,
	w108_0,w108_1,w108_2,w108_3,w108_4,w108_5,w108_6,w108_7,w108_8,w108_9,w108_10,w108_11,w108_12,w108_13,w108_14,w108_15,w108_16,
		w108_17,w108_18,w108_19,w108_20,w108_21,w108_22,w108_23,w108_24,w108_25,w108_26,w108_27,w108_28,w108_29,w108_30,w108_31,w108_32,
		w108_33,w108_34,w108_35,w108_36,w108_37,w108_38,w108_39,w108_40,w108_41,w108_42,w108_43,w108_44,w108_45,w108_46,w108_47,w108_48,
		w108_49,w108_50,w108_51,w108_52,w108_53,w108_54,w108_55,w108_56,w108_57,w108_58,w108_59,w108_60,w108_61,w108_62,w108_63,w108_64,
		w108_65,w108_66,w108_67,w108_68,w108_69,w108_70,w108_71,w108_72,w108_73,w108_74,w108_75,w108_76,w108_77,w108_78,w108_79,w108_80,
		w108_81,w108_82,w108_83,w108_84,w108_85,w108_86,w108_87,w108_88,w108_89,w108_90,w108_91,w108_92,w108_93,w108_94,w108_95,w108_96,
		w108_97,w108_98,w108_99,w108_100,w108_101,w108_102,w108_103,w108_104,w108_105,w108_106,w108_107,w108_108,w108_109,w108_110,w108_111,w108_112,
		w108_113,w108_114,w108_115,w108_116,w108_117,w108_118,w108_119,w108_120,w108_121,w108_122,w108_123,w108_124,w108_125,w108_126,
	w109_0,w109_1,w109_2,w109_3,w109_4,w109_5,w109_6,w109_7,w109_8,w109_9,w109_10,w109_11,w109_12,w109_13,w109_14,w109_15,w109_16,
		w109_17,w109_18,w109_19,w109_20,w109_21,w109_22,w109_23,w109_24,w109_25,w109_26,w109_27,w109_28,w109_29,w109_30,w109_31,w109_32,
		w109_33,w109_34,w109_35,w109_36,w109_37,w109_38,w109_39,w109_40,w109_41,w109_42,w109_43,w109_44,w109_45,w109_46,w109_47,w109_48,
		w109_49,w109_50,w109_51,w109_52,w109_53,w109_54,w109_55,w109_56,w109_57,w109_58,w109_59,w109_60,w109_61,w109_62,w109_63,w109_64,
		w109_65,w109_66,w109_67,w109_68,w109_69,w109_70,w109_71,w109_72,w109_73,w109_74,w109_75,w109_76,w109_77,w109_78,w109_79,w109_80,
		w109_81,w109_82,w109_83,w109_84,w109_85,w109_86,w109_87,w109_88,w109_89,w109_90,w109_91,w109_92,w109_93,w109_94,w109_95,w109_96,
		w109_97,w109_98,w109_99,w109_100,w109_101,w109_102,w109_103,w109_104,w109_105,w109_106,w109_107,w109_108,w109_109,w109_110,w109_111,w109_112,
		w109_113,w109_114,w109_115,w109_116,w109_117,w109_118,w109_119,w109_120,w109_121,w109_122,w109_123,w109_124,w109_125,w109_126,
	w110_0,w110_1,w110_2,w110_3,w110_4,w110_5,w110_6,w110_7,w110_8,w110_9,w110_10,w110_11,w110_12,w110_13,w110_14,w110_15,w110_16,
		w110_17,w110_18,w110_19,w110_20,w110_21,w110_22,w110_23,w110_24,w110_25,w110_26,w110_27,w110_28,w110_29,w110_30,w110_31,w110_32,
		w110_33,w110_34,w110_35,w110_36,w110_37,w110_38,w110_39,w110_40,w110_41,w110_42,w110_43,w110_44,w110_45,w110_46,w110_47,w110_48,
		w110_49,w110_50,w110_51,w110_52,w110_53,w110_54,w110_55,w110_56,w110_57,w110_58,w110_59,w110_60,w110_61,w110_62,w110_63,w110_64,
		w110_65,w110_66,w110_67,w110_68,w110_69,w110_70,w110_71,w110_72,w110_73,w110_74,w110_75,w110_76,w110_77,w110_78,w110_79,w110_80,
		w110_81,w110_82,w110_83,w110_84,w110_85,w110_86,w110_87,w110_88,w110_89,w110_90,w110_91,w110_92,w110_93,w110_94,w110_95,w110_96,
		w110_97,w110_98,w110_99,w110_100,w110_101,w110_102,w110_103,w110_104,w110_105,w110_106,w110_107,w110_108,w110_109,w110_110,w110_111,w110_112,
		w110_113,w110_114,w110_115,w110_116,w110_117,w110_118,w110_119,w110_120,w110_121,w110_122,w110_123,w110_124,w110_125,w110_126,
	w111_0,w111_1,w111_2,w111_3,w111_4,w111_5,w111_6,w111_7,w111_8,w111_9,w111_10,w111_11,w111_12,w111_13,w111_14,w111_15,w111_16,
		w111_17,w111_18,w111_19,w111_20,w111_21,w111_22,w111_23,w111_24,w111_25,w111_26,w111_27,w111_28,w111_29,w111_30,w111_31,w111_32,
		w111_33,w111_34,w111_35,w111_36,w111_37,w111_38,w111_39,w111_40,w111_41,w111_42,w111_43,w111_44,w111_45,w111_46,w111_47,w111_48,
		w111_49,w111_50,w111_51,w111_52,w111_53,w111_54,w111_55,w111_56,w111_57,w111_58,w111_59,w111_60,w111_61,w111_62,w111_63,w111_64,
		w111_65,w111_66,w111_67,w111_68,w111_69,w111_70,w111_71,w111_72,w111_73,w111_74,w111_75,w111_76,w111_77,w111_78,w111_79,w111_80,
		w111_81,w111_82,w111_83,w111_84,w111_85,w111_86,w111_87,w111_88,w111_89,w111_90,w111_91,w111_92,w111_93,w111_94,w111_95,w111_96,
		w111_97,w111_98,w111_99,w111_100,w111_101,w111_102,w111_103,w111_104,w111_105,w111_106,w111_107,w111_108,w111_109,w111_110,w111_111,w111_112,
		w111_113,w111_114,w111_115,w111_116,w111_117,w111_118,w111_119,w111_120,w111_121,w111_122,w111_123,w111_124,w111_125,w111_126,
	w112_0,w112_1,w112_2,w112_3,w112_4,w112_5,w112_6,w112_7,w112_8,w112_9,w112_10,w112_11,w112_12,w112_13,w112_14,w112_15,w112_16,
		w112_17,w112_18,w112_19,w112_20,w112_21,w112_22,w112_23,w112_24,w112_25,w112_26,w112_27,w112_28,w112_29,w112_30,w112_31,w112_32,
		w112_33,w112_34,w112_35,w112_36,w112_37,w112_38,w112_39,w112_40,w112_41,w112_42,w112_43,w112_44,w112_45,w112_46,w112_47,w112_48,
		w112_49,w112_50,w112_51,w112_52,w112_53,w112_54,w112_55,w112_56,w112_57,w112_58,w112_59,w112_60,w112_61,w112_62,w112_63,w112_64,
		w112_65,w112_66,w112_67,w112_68,w112_69,w112_70,w112_71,w112_72,w112_73,w112_74,w112_75,w112_76,w112_77,w112_78,w112_79,w112_80,
		w112_81,w112_82,w112_83,w112_84,w112_85,w112_86,w112_87,w112_88,w112_89,w112_90,w112_91,w112_92,w112_93,w112_94,w112_95,w112_96,
		w112_97,w112_98,w112_99,w112_100,w112_101,w112_102,w112_103,w112_104,w112_105,w112_106,w112_107,w112_108,w112_109,w112_110,w112_111,w112_112,
		w112_113,w112_114,w112_115,w112_116,w112_117,w112_118,w112_119,w112_120,w112_121,w112_122,w112_123,w112_124,w112_125,w112_126,
	w113_0,w113_1,w113_2,w113_3,w113_4,w113_5,w113_6,w113_7,w113_8,w113_9,w113_10,w113_11,w113_12,w113_13,w113_14,w113_15,w113_16,
		w113_17,w113_18,w113_19,w113_20,w113_21,w113_22,w113_23,w113_24,w113_25,w113_26,w113_27,w113_28,w113_29,w113_30,w113_31,w113_32,
		w113_33,w113_34,w113_35,w113_36,w113_37,w113_38,w113_39,w113_40,w113_41,w113_42,w113_43,w113_44,w113_45,w113_46,w113_47,w113_48,
		w113_49,w113_50,w113_51,w113_52,w113_53,w113_54,w113_55,w113_56,w113_57,w113_58,w113_59,w113_60,w113_61,w113_62,w113_63,w113_64,
		w113_65,w113_66,w113_67,w113_68,w113_69,w113_70,w113_71,w113_72,w113_73,w113_74,w113_75,w113_76,w113_77,w113_78,w113_79,w113_80,
		w113_81,w113_82,w113_83,w113_84,w113_85,w113_86,w113_87,w113_88,w113_89,w113_90,w113_91,w113_92,w113_93,w113_94,w113_95,w113_96,
		w113_97,w113_98,w113_99,w113_100,w113_101,w113_102,w113_103,w113_104,w113_105,w113_106,w113_107,w113_108,w113_109,w113_110,w113_111,w113_112,
		w113_113,w113_114,w113_115,w113_116,w113_117,w113_118,w113_119,w113_120,w113_121,w113_122,w113_123,w113_124,w113_125,w113_126,
	w114_0,w114_1,w114_2,w114_3,w114_4,w114_5,w114_6,w114_7,w114_8,w114_9,w114_10,w114_11,w114_12,w114_13,w114_14,w114_15,w114_16,
		w114_17,w114_18,w114_19,w114_20,w114_21,w114_22,w114_23,w114_24,w114_25,w114_26,w114_27,w114_28,w114_29,w114_30,w114_31,w114_32,
		w114_33,w114_34,w114_35,w114_36,w114_37,w114_38,w114_39,w114_40,w114_41,w114_42,w114_43,w114_44,w114_45,w114_46,w114_47,w114_48,
		w114_49,w114_50,w114_51,w114_52,w114_53,w114_54,w114_55,w114_56,w114_57,w114_58,w114_59,w114_60,w114_61,w114_62,w114_63,w114_64,
		w114_65,w114_66,w114_67,w114_68,w114_69,w114_70,w114_71,w114_72,w114_73,w114_74,w114_75,w114_76,w114_77,w114_78,w114_79,w114_80,
		w114_81,w114_82,w114_83,w114_84,w114_85,w114_86,w114_87,w114_88,w114_89,w114_90,w114_91,w114_92,w114_93,w114_94,w114_95,w114_96,
		w114_97,w114_98,w114_99,w114_100,w114_101,w114_102,w114_103,w114_104,w114_105,w114_106,w114_107,w114_108,w114_109,w114_110,w114_111,w114_112,
		w114_113,w114_114,w114_115,w114_116,w114_117,w114_118,w114_119,w114_120,w114_121,w114_122,w114_123,w114_124,w114_125,w114_126,
	w115_0,w115_1,w115_2,w115_3,w115_4,w115_5,w115_6,w115_7,w115_8,w115_9,w115_10,w115_11,w115_12,w115_13,w115_14,w115_15,w115_16,
		w115_17,w115_18,w115_19,w115_20,w115_21,w115_22,w115_23,w115_24,w115_25,w115_26,w115_27,w115_28,w115_29,w115_30,w115_31,w115_32,
		w115_33,w115_34,w115_35,w115_36,w115_37,w115_38,w115_39,w115_40,w115_41,w115_42,w115_43,w115_44,w115_45,w115_46,w115_47,w115_48,
		w115_49,w115_50,w115_51,w115_52,w115_53,w115_54,w115_55,w115_56,w115_57,w115_58,w115_59,w115_60,w115_61,w115_62,w115_63,w115_64,
		w115_65,w115_66,w115_67,w115_68,w115_69,w115_70,w115_71,w115_72,w115_73,w115_74,w115_75,w115_76,w115_77,w115_78,w115_79,w115_80,
		w115_81,w115_82,w115_83,w115_84,w115_85,w115_86,w115_87,w115_88,w115_89,w115_90,w115_91,w115_92,w115_93,w115_94,w115_95,w115_96,
		w115_97,w115_98,w115_99,w115_100,w115_101,w115_102,w115_103,w115_104,w115_105,w115_106,w115_107,w115_108,w115_109,w115_110,w115_111,w115_112,
		w115_113,w115_114,w115_115,w115_116,w115_117,w115_118,w115_119,w115_120,w115_121,w115_122,w115_123,w115_124,w115_125,w115_126,
	w116_0,w116_1,w116_2,w116_3,w116_4,w116_5,w116_6,w116_7,w116_8,w116_9,w116_10,w116_11,w116_12,w116_13,w116_14,w116_15,w116_16,
		w116_17,w116_18,w116_19,w116_20,w116_21,w116_22,w116_23,w116_24,w116_25,w116_26,w116_27,w116_28,w116_29,w116_30,w116_31,w116_32,
		w116_33,w116_34,w116_35,w116_36,w116_37,w116_38,w116_39,w116_40,w116_41,w116_42,w116_43,w116_44,w116_45,w116_46,w116_47,w116_48,
		w116_49,w116_50,w116_51,w116_52,w116_53,w116_54,w116_55,w116_56,w116_57,w116_58,w116_59,w116_60,w116_61,w116_62,w116_63,w116_64,
		w116_65,w116_66,w116_67,w116_68,w116_69,w116_70,w116_71,w116_72,w116_73,w116_74,w116_75,w116_76,w116_77,w116_78,w116_79,w116_80,
		w116_81,w116_82,w116_83,w116_84,w116_85,w116_86,w116_87,w116_88,w116_89,w116_90,w116_91,w116_92,w116_93,w116_94,w116_95,w116_96,
		w116_97,w116_98,w116_99,w116_100,w116_101,w116_102,w116_103,w116_104,w116_105,w116_106,w116_107,w116_108,w116_109,w116_110,w116_111,w116_112,
		w116_113,w116_114,w116_115,w116_116,w116_117,w116_118,w116_119,w116_120,w116_121,w116_122,w116_123,w116_124,w116_125,w116_126,
	w117_0,w117_1,w117_2,w117_3,w117_4,w117_5,w117_6,w117_7,w117_8,w117_9,w117_10,w117_11,w117_12,w117_13,w117_14,w117_15,w117_16,
		w117_17,w117_18,w117_19,w117_20,w117_21,w117_22,w117_23,w117_24,w117_25,w117_26,w117_27,w117_28,w117_29,w117_30,w117_31,w117_32,
		w117_33,w117_34,w117_35,w117_36,w117_37,w117_38,w117_39,w117_40,w117_41,w117_42,w117_43,w117_44,w117_45,w117_46,w117_47,w117_48,
		w117_49,w117_50,w117_51,w117_52,w117_53,w117_54,w117_55,w117_56,w117_57,w117_58,w117_59,w117_60,w117_61,w117_62,w117_63,w117_64,
		w117_65,w117_66,w117_67,w117_68,w117_69,w117_70,w117_71,w117_72,w117_73,w117_74,w117_75,w117_76,w117_77,w117_78,w117_79,w117_80,
		w117_81,w117_82,w117_83,w117_84,w117_85,w117_86,w117_87,w117_88,w117_89,w117_90,w117_91,w117_92,w117_93,w117_94,w117_95,w117_96,
		w117_97,w117_98,w117_99,w117_100,w117_101,w117_102,w117_103,w117_104,w117_105,w117_106,w117_107,w117_108,w117_109,w117_110,w117_111,w117_112,
		w117_113,w117_114,w117_115,w117_116,w117_117,w117_118,w117_119,w117_120,w117_121,w117_122,w117_123,w117_124,w117_125,w117_126,
	w118_0,w118_1,w118_2,w118_3,w118_4,w118_5,w118_6,w118_7,w118_8,w118_9,w118_10,w118_11,w118_12,w118_13,w118_14,w118_15,w118_16,
		w118_17,w118_18,w118_19,w118_20,w118_21,w118_22,w118_23,w118_24,w118_25,w118_26,w118_27,w118_28,w118_29,w118_30,w118_31,w118_32,
		w118_33,w118_34,w118_35,w118_36,w118_37,w118_38,w118_39,w118_40,w118_41,w118_42,w118_43,w118_44,w118_45,w118_46,w118_47,w118_48,
		w118_49,w118_50,w118_51,w118_52,w118_53,w118_54,w118_55,w118_56,w118_57,w118_58,w118_59,w118_60,w118_61,w118_62,w118_63,w118_64,
		w118_65,w118_66,w118_67,w118_68,w118_69,w118_70,w118_71,w118_72,w118_73,w118_74,w118_75,w118_76,w118_77,w118_78,w118_79,w118_80,
		w118_81,w118_82,w118_83,w118_84,w118_85,w118_86,w118_87,w118_88,w118_89,w118_90,w118_91,w118_92,w118_93,w118_94,w118_95,w118_96,
		w118_97,w118_98,w118_99,w118_100,w118_101,w118_102,w118_103,w118_104,w118_105,w118_106,w118_107,w118_108,w118_109,w118_110,w118_111,w118_112,
		w118_113,w118_114,w118_115,w118_116,w118_117,w118_118,w118_119,w118_120,w118_121,w118_122,w118_123,w118_124,w118_125,w118_126,
	w119_0,w119_1,w119_2,w119_3,w119_4,w119_5,w119_6,w119_7,w119_8,w119_9,w119_10,w119_11,w119_12,w119_13,w119_14,w119_15,w119_16,
		w119_17,w119_18,w119_19,w119_20,w119_21,w119_22,w119_23,w119_24,w119_25,w119_26,w119_27,w119_28,w119_29,w119_30,w119_31,w119_32,
		w119_33,w119_34,w119_35,w119_36,w119_37,w119_38,w119_39,w119_40,w119_41,w119_42,w119_43,w119_44,w119_45,w119_46,w119_47,w119_48,
		w119_49,w119_50,w119_51,w119_52,w119_53,w119_54,w119_55,w119_56,w119_57,w119_58,w119_59,w119_60,w119_61,w119_62,w119_63,w119_64,
		w119_65,w119_66,w119_67,w119_68,w119_69,w119_70,w119_71,w119_72,w119_73,w119_74,w119_75,w119_76,w119_77,w119_78,w119_79,w119_80,
		w119_81,w119_82,w119_83,w119_84,w119_85,w119_86,w119_87,w119_88,w119_89,w119_90,w119_91,w119_92,w119_93,w119_94,w119_95,w119_96,
		w119_97,w119_98,w119_99,w119_100,w119_101,w119_102,w119_103,w119_104,w119_105,w119_106,w119_107,w119_108,w119_109,w119_110,w119_111,w119_112,
		w119_113,w119_114,w119_115,w119_116,w119_117,w119_118,w119_119,w119_120,w119_121,w119_122,w119_123,w119_124,w119_125,w119_126,
	w120_0,w120_1,w120_2,w120_3,w120_4,w120_5,w120_6,w120_7,w120_8,w120_9,w120_10,w120_11,w120_12,w120_13,w120_14,w120_15,w120_16,
		w120_17,w120_18,w120_19,w120_20,w120_21,w120_22,w120_23,w120_24,w120_25,w120_26,w120_27,w120_28,w120_29,w120_30,w120_31,w120_32,
		w120_33,w120_34,w120_35,w120_36,w120_37,w120_38,w120_39,w120_40,w120_41,w120_42,w120_43,w120_44,w120_45,w120_46,w120_47,w120_48,
		w120_49,w120_50,w120_51,w120_52,w120_53,w120_54,w120_55,w120_56,w120_57,w120_58,w120_59,w120_60,w120_61,w120_62,w120_63,w120_64,
		w120_65,w120_66,w120_67,w120_68,w120_69,w120_70,w120_71,w120_72,w120_73,w120_74,w120_75,w120_76,w120_77,w120_78,w120_79,w120_80,
		w120_81,w120_82,w120_83,w120_84,w120_85,w120_86,w120_87,w120_88,w120_89,w120_90,w120_91,w120_92,w120_93,w120_94,w120_95,w120_96,
		w120_97,w120_98,w120_99,w120_100,w120_101,w120_102,w120_103,w120_104,w120_105,w120_106,w120_107,w120_108,w120_109,w120_110,w120_111,w120_112,
		w120_113,w120_114,w120_115,w120_116,w120_117,w120_118,w120_119,w120_120,w120_121,w120_122,w120_123,w120_124,w120_125,w120_126,
	w121_0,w121_1,w121_2,w121_3,w121_4,w121_5,w121_6,w121_7,w121_8,w121_9,w121_10,w121_11,w121_12,w121_13,w121_14,w121_15,w121_16,
		w121_17,w121_18,w121_19,w121_20,w121_21,w121_22,w121_23,w121_24,w121_25,w121_26,w121_27,w121_28,w121_29,w121_30,w121_31,w121_32,
		w121_33,w121_34,w121_35,w121_36,w121_37,w121_38,w121_39,w121_40,w121_41,w121_42,w121_43,w121_44,w121_45,w121_46,w121_47,w121_48,
		w121_49,w121_50,w121_51,w121_52,w121_53,w121_54,w121_55,w121_56,w121_57,w121_58,w121_59,w121_60,w121_61,w121_62,w121_63,w121_64,
		w121_65,w121_66,w121_67,w121_68,w121_69,w121_70,w121_71,w121_72,w121_73,w121_74,w121_75,w121_76,w121_77,w121_78,w121_79,w121_80,
		w121_81,w121_82,w121_83,w121_84,w121_85,w121_86,w121_87,w121_88,w121_89,w121_90,w121_91,w121_92,w121_93,w121_94,w121_95,w121_96,
		w121_97,w121_98,w121_99,w121_100,w121_101,w121_102,w121_103,w121_104,w121_105,w121_106,w121_107,w121_108,w121_109,w121_110,w121_111,w121_112,
		w121_113,w121_114,w121_115,w121_116,w121_117,w121_118,w121_119,w121_120,w121_121,w121_122,w121_123,w121_124,w121_125,w121_126,
	w122_0,w122_1,w122_2,w122_3,w122_4,w122_5,w122_6,w122_7,w122_8,w122_9,w122_10,w122_11,w122_12,w122_13,w122_14,w122_15,w122_16,
		w122_17,w122_18,w122_19,w122_20,w122_21,w122_22,w122_23,w122_24,w122_25,w122_26,w122_27,w122_28,w122_29,w122_30,w122_31,w122_32,
		w122_33,w122_34,w122_35,w122_36,w122_37,w122_38,w122_39,w122_40,w122_41,w122_42,w122_43,w122_44,w122_45,w122_46,w122_47,w122_48,
		w122_49,w122_50,w122_51,w122_52,w122_53,w122_54,w122_55,w122_56,w122_57,w122_58,w122_59,w122_60,w122_61,w122_62,w122_63,w122_64,
		w122_65,w122_66,w122_67,w122_68,w122_69,w122_70,w122_71,w122_72,w122_73,w122_74,w122_75,w122_76,w122_77,w122_78,w122_79,w122_80,
		w122_81,w122_82,w122_83,w122_84,w122_85,w122_86,w122_87,w122_88,w122_89,w122_90,w122_91,w122_92,w122_93,w122_94,w122_95,w122_96,
		w122_97,w122_98,w122_99,w122_100,w122_101,w122_102,w122_103,w122_104,w122_105,w122_106,w122_107,w122_108,w122_109,w122_110,w122_111,w122_112,
		w122_113,w122_114,w122_115,w122_116,w122_117,w122_118,w122_119,w122_120,w122_121,w122_122,w122_123,w122_124,w122_125,w122_126,
	w123_0,w123_1,w123_2,w123_3,w123_4,w123_5,w123_6,w123_7,w123_8,w123_9,w123_10,w123_11,w123_12,w123_13,w123_14,w123_15,w123_16,
		w123_17,w123_18,w123_19,w123_20,w123_21,w123_22,w123_23,w123_24,w123_25,w123_26,w123_27,w123_28,w123_29,w123_30,w123_31,w123_32,
		w123_33,w123_34,w123_35,w123_36,w123_37,w123_38,w123_39,w123_40,w123_41,w123_42,w123_43,w123_44,w123_45,w123_46,w123_47,w123_48,
		w123_49,w123_50,w123_51,w123_52,w123_53,w123_54,w123_55,w123_56,w123_57,w123_58,w123_59,w123_60,w123_61,w123_62,w123_63,w123_64,
		w123_65,w123_66,w123_67,w123_68,w123_69,w123_70,w123_71,w123_72,w123_73,w123_74,w123_75,w123_76,w123_77,w123_78,w123_79,w123_80,
		w123_81,w123_82,w123_83,w123_84,w123_85,w123_86,w123_87,w123_88,w123_89,w123_90,w123_91,w123_92,w123_93,w123_94,w123_95,w123_96,
		w123_97,w123_98,w123_99,w123_100,w123_101,w123_102,w123_103,w123_104,w123_105,w123_106,w123_107,w123_108,w123_109,w123_110,w123_111,w123_112,
		w123_113,w123_114,w123_115,w123_116,w123_117,w123_118,w123_119,w123_120,w123_121,w123_122,w123_123,w123_124,w123_125,w123_126,
	w124_0,w124_1,w124_2,w124_3,w124_4,w124_5,w124_6,w124_7,w124_8,w124_9,w124_10,w124_11,w124_12,w124_13,w124_14,w124_15,w124_16,
		w124_17,w124_18,w124_19,w124_20,w124_21,w124_22,w124_23,w124_24,w124_25,w124_26,w124_27,w124_28,w124_29,w124_30,w124_31,w124_32,
		w124_33,w124_34,w124_35,w124_36,w124_37,w124_38,w124_39,w124_40,w124_41,w124_42,w124_43,w124_44,w124_45,w124_46,w124_47,w124_48,
		w124_49,w124_50,w124_51,w124_52,w124_53,w124_54,w124_55,w124_56,w124_57,w124_58,w124_59,w124_60,w124_61,w124_62,w124_63,w124_64,
		w124_65,w124_66,w124_67,w124_68,w124_69,w124_70,w124_71,w124_72,w124_73,w124_74,w124_75,w124_76,w124_77,w124_78,w124_79,w124_80,
		w124_81,w124_82,w124_83,w124_84,w124_85,w124_86,w124_87,w124_88,w124_89,w124_90,w124_91,w124_92,w124_93,w124_94,w124_95,w124_96,
		w124_97,w124_98,w124_99,w124_100,w124_101,w124_102,w124_103,w124_104,w124_105,w124_106,w124_107,w124_108,w124_109,w124_110,w124_111,w124_112,
		w124_113,w124_114,w124_115,w124_116,w124_117,w124_118,w124_119,w124_120,w124_121,w124_122,w124_123,w124_124,w124_125,w124_126,
	w125_0,w125_1,w125_2,w125_3,w125_4,w125_5,w125_6,w125_7,w125_8,w125_9,w125_10,w125_11,w125_12,w125_13,w125_14,w125_15,w125_16,
		w125_17,w125_18,w125_19,w125_20,w125_21,w125_22,w125_23,w125_24,w125_25,w125_26,w125_27,w125_28,w125_29,w125_30,w125_31,w125_32,
		w125_33,w125_34,w125_35,w125_36,w125_37,w125_38,w125_39,w125_40,w125_41,w125_42,w125_43,w125_44,w125_45,w125_46,w125_47,w125_48,
		w125_49,w125_50,w125_51,w125_52,w125_53,w125_54,w125_55,w125_56,w125_57,w125_58,w125_59,w125_60,w125_61,w125_62,w125_63,w125_64,
		w125_65,w125_66,w125_67,w125_68,w125_69,w125_70,w125_71,w125_72,w125_73,w125_74,w125_75,w125_76,w125_77,w125_78,w125_79,w125_80,
		w125_81,w125_82,w125_83,w125_84,w125_85,w125_86,w125_87,w125_88,w125_89,w125_90,w125_91,w125_92,w125_93,w125_94,w125_95,w125_96,
		w125_97,w125_98,w125_99,w125_100,w125_101,w125_102,w125_103,w125_104,w125_105,w125_106,w125_107,w125_108,w125_109,w125_110,w125_111,w125_112,
		w125_113,w125_114,w125_115,w125_116,w125_117,w125_118,w125_119,w125_120,w125_121,w125_122,w125_123,w125_124,w125_125,w125_126,
	w126_0,w126_1,w126_2,w126_3,w126_4,w126_5,w126_6,w126_7,w126_8,w126_9,w126_10,w126_11,w126_12,w126_13,w126_14,w126_15,w126_16,
		w126_17,w126_18,w126_19,w126_20,w126_21,w126_22,w126_23,w126_24,w126_25,w126_26,w126_27,w126_28,w126_29,w126_30,w126_31,w126_32,
		w126_33,w126_34,w126_35,w126_36,w126_37,w126_38,w126_39,w126_40,w126_41,w126_42,w126_43,w126_44,w126_45,w126_46,w126_47,w126_48,
		w126_49,w126_50,w126_51,w126_52,w126_53,w126_54,w126_55,w126_56,w126_57,w126_58,w126_59,w126_60,w126_61,w126_62,w126_63,w126_64,
		w126_65,w126_66,w126_67,w126_68,w126_69,w126_70,w126_71,w126_72,w126_73,w126_74,w126_75,w126_76,w126_77,w126_78,w126_79,w126_80,
		w126_81,w126_82,w126_83,w126_84,w126_85,w126_86,w126_87,w126_88,w126_89,w126_90,w126_91,w126_92,w126_93,w126_94,w126_95,w126_96,
		w126_97,w126_98,w126_99,w126_100,w126_101,w126_102,w126_103,w126_104,w126_105,w126_106,w126_107,w126_108,w126_109,w126_110,w126_111,w126_112,
		w126_113,w126_114,w126_115,w126_116,w126_117,w126_118,w126_119,w126_120,w126_121,w126_122,w126_123,w126_124,w126_125,w126_126,
	w127_0,w127_1,w127_2,w127_3,w127_4,w127_5,w127_6,w127_7,w127_8,w127_9,w127_10,w127_11,w127_12,w127_13,w127_14,w127_15,w127_16,
		w127_17,w127_18,w127_19,w127_20,w127_21,w127_22,w127_23,w127_24,w127_25,w127_26,w127_27,w127_28,w127_29,w127_30,w127_31,w127_32,
		w127_33,w127_34,w127_35,w127_36,w127_37,w127_38,w127_39,w127_40,w127_41,w127_42,w127_43,w127_44,w127_45,w127_46,w127_47,w127_48,
		w127_49,w127_50,w127_51,w127_52,w127_53,w127_54,w127_55,w127_56,w127_57,w127_58,w127_59,w127_60,w127_61,w127_62,w127_63,w127_64,
		w127_65,w127_66,w127_67,w127_68,w127_69,w127_70,w127_71,w127_72,w127_73,w127_74,w127_75,w127_76,w127_77,w127_78,w127_79,w127_80,
		w127_81,w127_82,w127_83,w127_84,w127_85,w127_86,w127_87,w127_88,w127_89,w127_90,w127_91,w127_92,w127_93,w127_94,w127_95,w127_96,
		w127_97,w127_98,w127_99,w127_100,w127_101,w127_102,w127_103,w127_104,w127_105,w127_106,w127_107,w127_108,w127_109,w127_110,w127_111,w127_112,
		w127_113,w127_114,w127_115,w127_116,w127_117,w127_118,w127_119,w127_120,w127_121,w127_122,w127_123,w127_124,w127_125,w127_126;
	

	wire [31:0] r0_0,r0_1,r0_2,r0_3,r0_4,r0_5,r0_6,r0_7,r0_8,r0_9,r0_10,r0_11,r0_12,r0_13,r0_14,r0_15,r0_16,
		r0_17,r0_18,r0_19,r0_20,r0_21,r0_22,r0_23,r0_24,r0_25,r0_26,r0_27,r0_28,r0_29,r0_30,r0_31,r0_32,
		r0_33,r0_34,r0_35,r0_36,r0_37,r0_38,r0_39,r0_40,r0_41,r0_42,r0_43,r0_44,r0_45,r0_46,r0_47,r0_48,
		r0_49,r0_50,r0_51,r0_52,r0_53,r0_54,r0_55,r0_56,r0_57,r0_58,r0_59,r0_60,r0_61,r0_62,r0_63,r0_64,
		r0_65,r0_66,r0_67,r0_68,r0_69,r0_70,r0_71,r0_72,r0_73,r0_74,r0_75,r0_76,r0_77,r0_78,r0_79,r0_80,
		r0_81,r0_82,r0_83,r0_84,r0_85,r0_86,r0_87,r0_88,r0_89,r0_90,r0_91,r0_92,r0_93,r0_94,r0_95,r0_96,
		r0_97,r0_98,r0_99,r0_100,r0_101,r0_102,r0_103,r0_104,r0_105,r0_106,r0_107,r0_108,r0_109,r0_110,r0_111,r0_112,
		r0_113,r0_114,r0_115,r0_116,r0_117,r0_118,r0_119,r0_120,r0_121,r0_122,r0_123,r0_124,r0_125,r0_126,
	r1_0,r1_1,r1_2,r1_3,r1_4,r1_5,r1_6,r1_7,r1_8,r1_9,r1_10,r1_11,r1_12,r1_13,r1_14,r1_15,r1_16,
		r1_17,r1_18,r1_19,r1_20,r1_21,r1_22,r1_23,r1_24,r1_25,r1_26,r1_27,r1_28,r1_29,r1_30,r1_31,r1_32,
		r1_33,r1_34,r1_35,r1_36,r1_37,r1_38,r1_39,r1_40,r1_41,r1_42,r1_43,r1_44,r1_45,r1_46,r1_47,r1_48,
		r1_49,r1_50,r1_51,r1_52,r1_53,r1_54,r1_55,r1_56,r1_57,r1_58,r1_59,r1_60,r1_61,r1_62,r1_63,r1_64,
		r1_65,r1_66,r1_67,r1_68,r1_69,r1_70,r1_71,r1_72,r1_73,r1_74,r1_75,r1_76,r1_77,r1_78,r1_79,r1_80,
		r1_81,r1_82,r1_83,r1_84,r1_85,r1_86,r1_87,r1_88,r1_89,r1_90,r1_91,r1_92,r1_93,r1_94,r1_95,r1_96,
		r1_97,r1_98,r1_99,r1_100,r1_101,r1_102,r1_103,r1_104,r1_105,r1_106,r1_107,r1_108,r1_109,r1_110,r1_111,r1_112,
		r1_113,r1_114,r1_115,r1_116,r1_117,r1_118,r1_119,r1_120,r1_121,r1_122,r1_123,r1_124,r1_125,r1_126,
	r2_0,r2_1,r2_2,r2_3,r2_4,r2_5,r2_6,r2_7,r2_8,r2_9,r2_10,r2_11,r2_12,r2_13,r2_14,r2_15,r2_16,
		r2_17,r2_18,r2_19,r2_20,r2_21,r2_22,r2_23,r2_24,r2_25,r2_26,r2_27,r2_28,r2_29,r2_30,r2_31,r2_32,
		r2_33,r2_34,r2_35,r2_36,r2_37,r2_38,r2_39,r2_40,r2_41,r2_42,r2_43,r2_44,r2_45,r2_46,r2_47,r2_48,
		r2_49,r2_50,r2_51,r2_52,r2_53,r2_54,r2_55,r2_56,r2_57,r2_58,r2_59,r2_60,r2_61,r2_62,r2_63,r2_64,
		r2_65,r2_66,r2_67,r2_68,r2_69,r2_70,r2_71,r2_72,r2_73,r2_74,r2_75,r2_76,r2_77,r2_78,r2_79,r2_80,
		r2_81,r2_82,r2_83,r2_84,r2_85,r2_86,r2_87,r2_88,r2_89,r2_90,r2_91,r2_92,r2_93,r2_94,r2_95,r2_96,
		r2_97,r2_98,r2_99,r2_100,r2_101,r2_102,r2_103,r2_104,r2_105,r2_106,r2_107,r2_108,r2_109,r2_110,r2_111,r2_112,
		r2_113,r2_114,r2_115,r2_116,r2_117,r2_118,r2_119,r2_120,r2_121,r2_122,r2_123,r2_124,r2_125,r2_126,
	r3_0,r3_1,r3_2,r3_3,r3_4,r3_5,r3_6,r3_7,r3_8,r3_9,r3_10,r3_11,r3_12,r3_13,r3_14,r3_15,r3_16,
		r3_17,r3_18,r3_19,r3_20,r3_21,r3_22,r3_23,r3_24,r3_25,r3_26,r3_27,r3_28,r3_29,r3_30,r3_31,r3_32,
		r3_33,r3_34,r3_35,r3_36,r3_37,r3_38,r3_39,r3_40,r3_41,r3_42,r3_43,r3_44,r3_45,r3_46,r3_47,r3_48,
		r3_49,r3_50,r3_51,r3_52,r3_53,r3_54,r3_55,r3_56,r3_57,r3_58,r3_59,r3_60,r3_61,r3_62,r3_63,r3_64,
		r3_65,r3_66,r3_67,r3_68,r3_69,r3_70,r3_71,r3_72,r3_73,r3_74,r3_75,r3_76,r3_77,r3_78,r3_79,r3_80,
		r3_81,r3_82,r3_83,r3_84,r3_85,r3_86,r3_87,r3_88,r3_89,r3_90,r3_91,r3_92,r3_93,r3_94,r3_95,r3_96,
		r3_97,r3_98,r3_99,r3_100,r3_101,r3_102,r3_103,r3_104,r3_105,r3_106,r3_107,r3_108,r3_109,r3_110,r3_111,r3_112,
		r3_113,r3_114,r3_115,r3_116,r3_117,r3_118,r3_119,r3_120,r3_121,r3_122,r3_123,r3_124,r3_125,r3_126,
	r4_0,r4_1,r4_2,r4_3,r4_4,r4_5,r4_6,r4_7,r4_8,r4_9,r4_10,r4_11,r4_12,r4_13,r4_14,r4_15,r4_16,
		r4_17,r4_18,r4_19,r4_20,r4_21,r4_22,r4_23,r4_24,r4_25,r4_26,r4_27,r4_28,r4_29,r4_30,r4_31,r4_32,
		r4_33,r4_34,r4_35,r4_36,r4_37,r4_38,r4_39,r4_40,r4_41,r4_42,r4_43,r4_44,r4_45,r4_46,r4_47,r4_48,
		r4_49,r4_50,r4_51,r4_52,r4_53,r4_54,r4_55,r4_56,r4_57,r4_58,r4_59,r4_60,r4_61,r4_62,r4_63,r4_64,
		r4_65,r4_66,r4_67,r4_68,r4_69,r4_70,r4_71,r4_72,r4_73,r4_74,r4_75,r4_76,r4_77,r4_78,r4_79,r4_80,
		r4_81,r4_82,r4_83,r4_84,r4_85,r4_86,r4_87,r4_88,r4_89,r4_90,r4_91,r4_92,r4_93,r4_94,r4_95,r4_96,
		r4_97,r4_98,r4_99,r4_100,r4_101,r4_102,r4_103,r4_104,r4_105,r4_106,r4_107,r4_108,r4_109,r4_110,r4_111,r4_112,
		r4_113,r4_114,r4_115,r4_116,r4_117,r4_118,r4_119,r4_120,r4_121,r4_122,r4_123,r4_124,r4_125,r4_126,
	r5_0,r5_1,r5_2,r5_3,r5_4,r5_5,r5_6,r5_7,r5_8,r5_9,r5_10,r5_11,r5_12,r5_13,r5_14,r5_15,r5_16,
		r5_17,r5_18,r5_19,r5_20,r5_21,r5_22,r5_23,r5_24,r5_25,r5_26,r5_27,r5_28,r5_29,r5_30,r5_31,r5_32,
		r5_33,r5_34,r5_35,r5_36,r5_37,r5_38,r5_39,r5_40,r5_41,r5_42,r5_43,r5_44,r5_45,r5_46,r5_47,r5_48,
		r5_49,r5_50,r5_51,r5_52,r5_53,r5_54,r5_55,r5_56,r5_57,r5_58,r5_59,r5_60,r5_61,r5_62,r5_63,r5_64,
		r5_65,r5_66,r5_67,r5_68,r5_69,r5_70,r5_71,r5_72,r5_73,r5_74,r5_75,r5_76,r5_77,r5_78,r5_79,r5_80,
		r5_81,r5_82,r5_83,r5_84,r5_85,r5_86,r5_87,r5_88,r5_89,r5_90,r5_91,r5_92,r5_93,r5_94,r5_95,r5_96,
		r5_97,r5_98,r5_99,r5_100,r5_101,r5_102,r5_103,r5_104,r5_105,r5_106,r5_107,r5_108,r5_109,r5_110,r5_111,r5_112,
		r5_113,r5_114,r5_115,r5_116,r5_117,r5_118,r5_119,r5_120,r5_121,r5_122,r5_123,r5_124,r5_125,r5_126,
	r6_0,r6_1,r6_2,r6_3,r6_4,r6_5,r6_6,r6_7,r6_8,r6_9,r6_10,r6_11,r6_12,r6_13,r6_14,r6_15,r6_16,
		r6_17,r6_18,r6_19,r6_20,r6_21,r6_22,r6_23,r6_24,r6_25,r6_26,r6_27,r6_28,r6_29,r6_30,r6_31,r6_32,
		r6_33,r6_34,r6_35,r6_36,r6_37,r6_38,r6_39,r6_40,r6_41,r6_42,r6_43,r6_44,r6_45,r6_46,r6_47,r6_48,
		r6_49,r6_50,r6_51,r6_52,r6_53,r6_54,r6_55,r6_56,r6_57,r6_58,r6_59,r6_60,r6_61,r6_62,r6_63,r6_64,
		r6_65,r6_66,r6_67,r6_68,r6_69,r6_70,r6_71,r6_72,r6_73,r6_74,r6_75,r6_76,r6_77,r6_78,r6_79,r6_80,
		r6_81,r6_82,r6_83,r6_84,r6_85,r6_86,r6_87,r6_88,r6_89,r6_90,r6_91,r6_92,r6_93,r6_94,r6_95,r6_96,
		r6_97,r6_98,r6_99,r6_100,r6_101,r6_102,r6_103,r6_104,r6_105,r6_106,r6_107,r6_108,r6_109,r6_110,r6_111,r6_112,
		r6_113,r6_114,r6_115,r6_116,r6_117,r6_118,r6_119,r6_120,r6_121,r6_122,r6_123,r6_124,r6_125,r6_126,
	r7_0,r7_1,r7_2,r7_3,r7_4,r7_5,r7_6,r7_7,r7_8,r7_9,r7_10,r7_11,r7_12,r7_13,r7_14,r7_15,r7_16,
		r7_17,r7_18,r7_19,r7_20,r7_21,r7_22,r7_23,r7_24,r7_25,r7_26,r7_27,r7_28,r7_29,r7_30,r7_31,r7_32,
		r7_33,r7_34,r7_35,r7_36,r7_37,r7_38,r7_39,r7_40,r7_41,r7_42,r7_43,r7_44,r7_45,r7_46,r7_47,r7_48,
		r7_49,r7_50,r7_51,r7_52,r7_53,r7_54,r7_55,r7_56,r7_57,r7_58,r7_59,r7_60,r7_61,r7_62,r7_63,r7_64,
		r7_65,r7_66,r7_67,r7_68,r7_69,r7_70,r7_71,r7_72,r7_73,r7_74,r7_75,r7_76,r7_77,r7_78,r7_79,r7_80,
		r7_81,r7_82,r7_83,r7_84,r7_85,r7_86,r7_87,r7_88,r7_89,r7_90,r7_91,r7_92,r7_93,r7_94,r7_95,r7_96,
		r7_97,r7_98,r7_99,r7_100,r7_101,r7_102,r7_103,r7_104,r7_105,r7_106,r7_107,r7_108,r7_109,r7_110,r7_111,r7_112,
		r7_113,r7_114,r7_115,r7_116,r7_117,r7_118,r7_119,r7_120,r7_121,r7_122,r7_123,r7_124,r7_125,r7_126,
	r8_0,r8_1,r8_2,r8_3,r8_4,r8_5,r8_6,r8_7,r8_8,r8_9,r8_10,r8_11,r8_12,r8_13,r8_14,r8_15,r8_16,
		r8_17,r8_18,r8_19,r8_20,r8_21,r8_22,r8_23,r8_24,r8_25,r8_26,r8_27,r8_28,r8_29,r8_30,r8_31,r8_32,
		r8_33,r8_34,r8_35,r8_36,r8_37,r8_38,r8_39,r8_40,r8_41,r8_42,r8_43,r8_44,r8_45,r8_46,r8_47,r8_48,
		r8_49,r8_50,r8_51,r8_52,r8_53,r8_54,r8_55,r8_56,r8_57,r8_58,r8_59,r8_60,r8_61,r8_62,r8_63,r8_64,
		r8_65,r8_66,r8_67,r8_68,r8_69,r8_70,r8_71,r8_72,r8_73,r8_74,r8_75,r8_76,r8_77,r8_78,r8_79,r8_80,
		r8_81,r8_82,r8_83,r8_84,r8_85,r8_86,r8_87,r8_88,r8_89,r8_90,r8_91,r8_92,r8_93,r8_94,r8_95,r8_96,
		r8_97,r8_98,r8_99,r8_100,r8_101,r8_102,r8_103,r8_104,r8_105,r8_106,r8_107,r8_108,r8_109,r8_110,r8_111,r8_112,
		r8_113,r8_114,r8_115,r8_116,r8_117,r8_118,r8_119,r8_120,r8_121,r8_122,r8_123,r8_124,r8_125,r8_126,
	r9_0,r9_1,r9_2,r9_3,r9_4,r9_5,r9_6,r9_7,r9_8,r9_9,r9_10,r9_11,r9_12,r9_13,r9_14,r9_15,r9_16,
		r9_17,r9_18,r9_19,r9_20,r9_21,r9_22,r9_23,r9_24,r9_25,r9_26,r9_27,r9_28,r9_29,r9_30,r9_31,r9_32,
		r9_33,r9_34,r9_35,r9_36,r9_37,r9_38,r9_39,r9_40,r9_41,r9_42,r9_43,r9_44,r9_45,r9_46,r9_47,r9_48,
		r9_49,r9_50,r9_51,r9_52,r9_53,r9_54,r9_55,r9_56,r9_57,r9_58,r9_59,r9_60,r9_61,r9_62,r9_63,r9_64,
		r9_65,r9_66,r9_67,r9_68,r9_69,r9_70,r9_71,r9_72,r9_73,r9_74,r9_75,r9_76,r9_77,r9_78,r9_79,r9_80,
		r9_81,r9_82,r9_83,r9_84,r9_85,r9_86,r9_87,r9_88,r9_89,r9_90,r9_91,r9_92,r9_93,r9_94,r9_95,r9_96,
		r9_97,r9_98,r9_99,r9_100,r9_101,r9_102,r9_103,r9_104,r9_105,r9_106,r9_107,r9_108,r9_109,r9_110,r9_111,r9_112,
		r9_113,r9_114,r9_115,r9_116,r9_117,r9_118,r9_119,r9_120,r9_121,r9_122,r9_123,r9_124,r9_125,r9_126,
	r10_0,r10_1,r10_2,r10_3,r10_4,r10_5,r10_6,r10_7,r10_8,r10_9,r10_10,r10_11,r10_12,r10_13,r10_14,r10_15,r10_16,
		r10_17,r10_18,r10_19,r10_20,r10_21,r10_22,r10_23,r10_24,r10_25,r10_26,r10_27,r10_28,r10_29,r10_30,r10_31,r10_32,
		r10_33,r10_34,r10_35,r10_36,r10_37,r10_38,r10_39,r10_40,r10_41,r10_42,r10_43,r10_44,r10_45,r10_46,r10_47,r10_48,
		r10_49,r10_50,r10_51,r10_52,r10_53,r10_54,r10_55,r10_56,r10_57,r10_58,r10_59,r10_60,r10_61,r10_62,r10_63,r10_64,
		r10_65,r10_66,r10_67,r10_68,r10_69,r10_70,r10_71,r10_72,r10_73,r10_74,r10_75,r10_76,r10_77,r10_78,r10_79,r10_80,
		r10_81,r10_82,r10_83,r10_84,r10_85,r10_86,r10_87,r10_88,r10_89,r10_90,r10_91,r10_92,r10_93,r10_94,r10_95,r10_96,
		r10_97,r10_98,r10_99,r10_100,r10_101,r10_102,r10_103,r10_104,r10_105,r10_106,r10_107,r10_108,r10_109,r10_110,r10_111,r10_112,
		r10_113,r10_114,r10_115,r10_116,r10_117,r10_118,r10_119,r10_120,r10_121,r10_122,r10_123,r10_124,r10_125,r10_126,
	r11_0,r11_1,r11_2,r11_3,r11_4,r11_5,r11_6,r11_7,r11_8,r11_9,r11_10,r11_11,r11_12,r11_13,r11_14,r11_15,r11_16,
		r11_17,r11_18,r11_19,r11_20,r11_21,r11_22,r11_23,r11_24,r11_25,r11_26,r11_27,r11_28,r11_29,r11_30,r11_31,r11_32,
		r11_33,r11_34,r11_35,r11_36,r11_37,r11_38,r11_39,r11_40,r11_41,r11_42,r11_43,r11_44,r11_45,r11_46,r11_47,r11_48,
		r11_49,r11_50,r11_51,r11_52,r11_53,r11_54,r11_55,r11_56,r11_57,r11_58,r11_59,r11_60,r11_61,r11_62,r11_63,r11_64,
		r11_65,r11_66,r11_67,r11_68,r11_69,r11_70,r11_71,r11_72,r11_73,r11_74,r11_75,r11_76,r11_77,r11_78,r11_79,r11_80,
		r11_81,r11_82,r11_83,r11_84,r11_85,r11_86,r11_87,r11_88,r11_89,r11_90,r11_91,r11_92,r11_93,r11_94,r11_95,r11_96,
		r11_97,r11_98,r11_99,r11_100,r11_101,r11_102,r11_103,r11_104,r11_105,r11_106,r11_107,r11_108,r11_109,r11_110,r11_111,r11_112,
		r11_113,r11_114,r11_115,r11_116,r11_117,r11_118,r11_119,r11_120,r11_121,r11_122,r11_123,r11_124,r11_125,r11_126,
	r12_0,r12_1,r12_2,r12_3,r12_4,r12_5,r12_6,r12_7,r12_8,r12_9,r12_10,r12_11,r12_12,r12_13,r12_14,r12_15,r12_16,
		r12_17,r12_18,r12_19,r12_20,r12_21,r12_22,r12_23,r12_24,r12_25,r12_26,r12_27,r12_28,r12_29,r12_30,r12_31,r12_32,
		r12_33,r12_34,r12_35,r12_36,r12_37,r12_38,r12_39,r12_40,r12_41,r12_42,r12_43,r12_44,r12_45,r12_46,r12_47,r12_48,
		r12_49,r12_50,r12_51,r12_52,r12_53,r12_54,r12_55,r12_56,r12_57,r12_58,r12_59,r12_60,r12_61,r12_62,r12_63,r12_64,
		r12_65,r12_66,r12_67,r12_68,r12_69,r12_70,r12_71,r12_72,r12_73,r12_74,r12_75,r12_76,r12_77,r12_78,r12_79,r12_80,
		r12_81,r12_82,r12_83,r12_84,r12_85,r12_86,r12_87,r12_88,r12_89,r12_90,r12_91,r12_92,r12_93,r12_94,r12_95,r12_96,
		r12_97,r12_98,r12_99,r12_100,r12_101,r12_102,r12_103,r12_104,r12_105,r12_106,r12_107,r12_108,r12_109,r12_110,r12_111,r12_112,
		r12_113,r12_114,r12_115,r12_116,r12_117,r12_118,r12_119,r12_120,r12_121,r12_122,r12_123,r12_124,r12_125,r12_126,
	r13_0,r13_1,r13_2,r13_3,r13_4,r13_5,r13_6,r13_7,r13_8,r13_9,r13_10,r13_11,r13_12,r13_13,r13_14,r13_15,r13_16,
		r13_17,r13_18,r13_19,r13_20,r13_21,r13_22,r13_23,r13_24,r13_25,r13_26,r13_27,r13_28,r13_29,r13_30,r13_31,r13_32,
		r13_33,r13_34,r13_35,r13_36,r13_37,r13_38,r13_39,r13_40,r13_41,r13_42,r13_43,r13_44,r13_45,r13_46,r13_47,r13_48,
		r13_49,r13_50,r13_51,r13_52,r13_53,r13_54,r13_55,r13_56,r13_57,r13_58,r13_59,r13_60,r13_61,r13_62,r13_63,r13_64,
		r13_65,r13_66,r13_67,r13_68,r13_69,r13_70,r13_71,r13_72,r13_73,r13_74,r13_75,r13_76,r13_77,r13_78,r13_79,r13_80,
		r13_81,r13_82,r13_83,r13_84,r13_85,r13_86,r13_87,r13_88,r13_89,r13_90,r13_91,r13_92,r13_93,r13_94,r13_95,r13_96,
		r13_97,r13_98,r13_99,r13_100,r13_101,r13_102,r13_103,r13_104,r13_105,r13_106,r13_107,r13_108,r13_109,r13_110,r13_111,r13_112,
		r13_113,r13_114,r13_115,r13_116,r13_117,r13_118,r13_119,r13_120,r13_121,r13_122,r13_123,r13_124,r13_125,r13_126,
	r14_0,r14_1,r14_2,r14_3,r14_4,r14_5,r14_6,r14_7,r14_8,r14_9,r14_10,r14_11,r14_12,r14_13,r14_14,r14_15,r14_16,
		r14_17,r14_18,r14_19,r14_20,r14_21,r14_22,r14_23,r14_24,r14_25,r14_26,r14_27,r14_28,r14_29,r14_30,r14_31,r14_32,
		r14_33,r14_34,r14_35,r14_36,r14_37,r14_38,r14_39,r14_40,r14_41,r14_42,r14_43,r14_44,r14_45,r14_46,r14_47,r14_48,
		r14_49,r14_50,r14_51,r14_52,r14_53,r14_54,r14_55,r14_56,r14_57,r14_58,r14_59,r14_60,r14_61,r14_62,r14_63,r14_64,
		r14_65,r14_66,r14_67,r14_68,r14_69,r14_70,r14_71,r14_72,r14_73,r14_74,r14_75,r14_76,r14_77,r14_78,r14_79,r14_80,
		r14_81,r14_82,r14_83,r14_84,r14_85,r14_86,r14_87,r14_88,r14_89,r14_90,r14_91,r14_92,r14_93,r14_94,r14_95,r14_96,
		r14_97,r14_98,r14_99,r14_100,r14_101,r14_102,r14_103,r14_104,r14_105,r14_106,r14_107,r14_108,r14_109,r14_110,r14_111,r14_112,
		r14_113,r14_114,r14_115,r14_116,r14_117,r14_118,r14_119,r14_120,r14_121,r14_122,r14_123,r14_124,r14_125,r14_126,
	r15_0,r15_1,r15_2,r15_3,r15_4,r15_5,r15_6,r15_7,r15_8,r15_9,r15_10,r15_11,r15_12,r15_13,r15_14,r15_15,r15_16,
		r15_17,r15_18,r15_19,r15_20,r15_21,r15_22,r15_23,r15_24,r15_25,r15_26,r15_27,r15_28,r15_29,r15_30,r15_31,r15_32,
		r15_33,r15_34,r15_35,r15_36,r15_37,r15_38,r15_39,r15_40,r15_41,r15_42,r15_43,r15_44,r15_45,r15_46,r15_47,r15_48,
		r15_49,r15_50,r15_51,r15_52,r15_53,r15_54,r15_55,r15_56,r15_57,r15_58,r15_59,r15_60,r15_61,r15_62,r15_63,r15_64,
		r15_65,r15_66,r15_67,r15_68,r15_69,r15_70,r15_71,r15_72,r15_73,r15_74,r15_75,r15_76,r15_77,r15_78,r15_79,r15_80,
		r15_81,r15_82,r15_83,r15_84,r15_85,r15_86,r15_87,r15_88,r15_89,r15_90,r15_91,r15_92,r15_93,r15_94,r15_95,r15_96,
		r15_97,r15_98,r15_99,r15_100,r15_101,r15_102,r15_103,r15_104,r15_105,r15_106,r15_107,r15_108,r15_109,r15_110,r15_111,r15_112,
		r15_113,r15_114,r15_115,r15_116,r15_117,r15_118,r15_119,r15_120,r15_121,r15_122,r15_123,r15_124,r15_125,r15_126,
	r16_0,r16_1,r16_2,r16_3,r16_4,r16_5,r16_6,r16_7,r16_8,r16_9,r16_10,r16_11,r16_12,r16_13,r16_14,r16_15,r16_16,
		r16_17,r16_18,r16_19,r16_20,r16_21,r16_22,r16_23,r16_24,r16_25,r16_26,r16_27,r16_28,r16_29,r16_30,r16_31,r16_32,
		r16_33,r16_34,r16_35,r16_36,r16_37,r16_38,r16_39,r16_40,r16_41,r16_42,r16_43,r16_44,r16_45,r16_46,r16_47,r16_48,
		r16_49,r16_50,r16_51,r16_52,r16_53,r16_54,r16_55,r16_56,r16_57,r16_58,r16_59,r16_60,r16_61,r16_62,r16_63,r16_64,
		r16_65,r16_66,r16_67,r16_68,r16_69,r16_70,r16_71,r16_72,r16_73,r16_74,r16_75,r16_76,r16_77,r16_78,r16_79,r16_80,
		r16_81,r16_82,r16_83,r16_84,r16_85,r16_86,r16_87,r16_88,r16_89,r16_90,r16_91,r16_92,r16_93,r16_94,r16_95,r16_96,
		r16_97,r16_98,r16_99,r16_100,r16_101,r16_102,r16_103,r16_104,r16_105,r16_106,r16_107,r16_108,r16_109,r16_110,r16_111,r16_112,
		r16_113,r16_114,r16_115,r16_116,r16_117,r16_118,r16_119,r16_120,r16_121,r16_122,r16_123,r16_124,r16_125,r16_126,
	r17_0,r17_1,r17_2,r17_3,r17_4,r17_5,r17_6,r17_7,r17_8,r17_9,r17_10,r17_11,r17_12,r17_13,r17_14,r17_15,r17_16,
		r17_17,r17_18,r17_19,r17_20,r17_21,r17_22,r17_23,r17_24,r17_25,r17_26,r17_27,r17_28,r17_29,r17_30,r17_31,r17_32,
		r17_33,r17_34,r17_35,r17_36,r17_37,r17_38,r17_39,r17_40,r17_41,r17_42,r17_43,r17_44,r17_45,r17_46,r17_47,r17_48,
		r17_49,r17_50,r17_51,r17_52,r17_53,r17_54,r17_55,r17_56,r17_57,r17_58,r17_59,r17_60,r17_61,r17_62,r17_63,r17_64,
		r17_65,r17_66,r17_67,r17_68,r17_69,r17_70,r17_71,r17_72,r17_73,r17_74,r17_75,r17_76,r17_77,r17_78,r17_79,r17_80,
		r17_81,r17_82,r17_83,r17_84,r17_85,r17_86,r17_87,r17_88,r17_89,r17_90,r17_91,r17_92,r17_93,r17_94,r17_95,r17_96,
		r17_97,r17_98,r17_99,r17_100,r17_101,r17_102,r17_103,r17_104,r17_105,r17_106,r17_107,r17_108,r17_109,r17_110,r17_111,r17_112,
		r17_113,r17_114,r17_115,r17_116,r17_117,r17_118,r17_119,r17_120,r17_121,r17_122,r17_123,r17_124,r17_125,r17_126,
	r18_0,r18_1,r18_2,r18_3,r18_4,r18_5,r18_6,r18_7,r18_8,r18_9,r18_10,r18_11,r18_12,r18_13,r18_14,r18_15,r18_16,
		r18_17,r18_18,r18_19,r18_20,r18_21,r18_22,r18_23,r18_24,r18_25,r18_26,r18_27,r18_28,r18_29,r18_30,r18_31,r18_32,
		r18_33,r18_34,r18_35,r18_36,r18_37,r18_38,r18_39,r18_40,r18_41,r18_42,r18_43,r18_44,r18_45,r18_46,r18_47,r18_48,
		r18_49,r18_50,r18_51,r18_52,r18_53,r18_54,r18_55,r18_56,r18_57,r18_58,r18_59,r18_60,r18_61,r18_62,r18_63,r18_64,
		r18_65,r18_66,r18_67,r18_68,r18_69,r18_70,r18_71,r18_72,r18_73,r18_74,r18_75,r18_76,r18_77,r18_78,r18_79,r18_80,
		r18_81,r18_82,r18_83,r18_84,r18_85,r18_86,r18_87,r18_88,r18_89,r18_90,r18_91,r18_92,r18_93,r18_94,r18_95,r18_96,
		r18_97,r18_98,r18_99,r18_100,r18_101,r18_102,r18_103,r18_104,r18_105,r18_106,r18_107,r18_108,r18_109,r18_110,r18_111,r18_112,
		r18_113,r18_114,r18_115,r18_116,r18_117,r18_118,r18_119,r18_120,r18_121,r18_122,r18_123,r18_124,r18_125,r18_126,
	r19_0,r19_1,r19_2,r19_3,r19_4,r19_5,r19_6,r19_7,r19_8,r19_9,r19_10,r19_11,r19_12,r19_13,r19_14,r19_15,r19_16,
		r19_17,r19_18,r19_19,r19_20,r19_21,r19_22,r19_23,r19_24,r19_25,r19_26,r19_27,r19_28,r19_29,r19_30,r19_31,r19_32,
		r19_33,r19_34,r19_35,r19_36,r19_37,r19_38,r19_39,r19_40,r19_41,r19_42,r19_43,r19_44,r19_45,r19_46,r19_47,r19_48,
		r19_49,r19_50,r19_51,r19_52,r19_53,r19_54,r19_55,r19_56,r19_57,r19_58,r19_59,r19_60,r19_61,r19_62,r19_63,r19_64,
		r19_65,r19_66,r19_67,r19_68,r19_69,r19_70,r19_71,r19_72,r19_73,r19_74,r19_75,r19_76,r19_77,r19_78,r19_79,r19_80,
		r19_81,r19_82,r19_83,r19_84,r19_85,r19_86,r19_87,r19_88,r19_89,r19_90,r19_91,r19_92,r19_93,r19_94,r19_95,r19_96,
		r19_97,r19_98,r19_99,r19_100,r19_101,r19_102,r19_103,r19_104,r19_105,r19_106,r19_107,r19_108,r19_109,r19_110,r19_111,r19_112,
		r19_113,r19_114,r19_115,r19_116,r19_117,r19_118,r19_119,r19_120,r19_121,r19_122,r19_123,r19_124,r19_125,r19_126,
	r20_0,r20_1,r20_2,r20_3,r20_4,r20_5,r20_6,r20_7,r20_8,r20_9,r20_10,r20_11,r20_12,r20_13,r20_14,r20_15,r20_16,
		r20_17,r20_18,r20_19,r20_20,r20_21,r20_22,r20_23,r20_24,r20_25,r20_26,r20_27,r20_28,r20_29,r20_30,r20_31,r20_32,
		r20_33,r20_34,r20_35,r20_36,r20_37,r20_38,r20_39,r20_40,r20_41,r20_42,r20_43,r20_44,r20_45,r20_46,r20_47,r20_48,
		r20_49,r20_50,r20_51,r20_52,r20_53,r20_54,r20_55,r20_56,r20_57,r20_58,r20_59,r20_60,r20_61,r20_62,r20_63,r20_64,
		r20_65,r20_66,r20_67,r20_68,r20_69,r20_70,r20_71,r20_72,r20_73,r20_74,r20_75,r20_76,r20_77,r20_78,r20_79,r20_80,
		r20_81,r20_82,r20_83,r20_84,r20_85,r20_86,r20_87,r20_88,r20_89,r20_90,r20_91,r20_92,r20_93,r20_94,r20_95,r20_96,
		r20_97,r20_98,r20_99,r20_100,r20_101,r20_102,r20_103,r20_104,r20_105,r20_106,r20_107,r20_108,r20_109,r20_110,r20_111,r20_112,
		r20_113,r20_114,r20_115,r20_116,r20_117,r20_118,r20_119,r20_120,r20_121,r20_122,r20_123,r20_124,r20_125,r20_126,
	r21_0,r21_1,r21_2,r21_3,r21_4,r21_5,r21_6,r21_7,r21_8,r21_9,r21_10,r21_11,r21_12,r21_13,r21_14,r21_15,r21_16,
		r21_17,r21_18,r21_19,r21_20,r21_21,r21_22,r21_23,r21_24,r21_25,r21_26,r21_27,r21_28,r21_29,r21_30,r21_31,r21_32,
		r21_33,r21_34,r21_35,r21_36,r21_37,r21_38,r21_39,r21_40,r21_41,r21_42,r21_43,r21_44,r21_45,r21_46,r21_47,r21_48,
		r21_49,r21_50,r21_51,r21_52,r21_53,r21_54,r21_55,r21_56,r21_57,r21_58,r21_59,r21_60,r21_61,r21_62,r21_63,r21_64,
		r21_65,r21_66,r21_67,r21_68,r21_69,r21_70,r21_71,r21_72,r21_73,r21_74,r21_75,r21_76,r21_77,r21_78,r21_79,r21_80,
		r21_81,r21_82,r21_83,r21_84,r21_85,r21_86,r21_87,r21_88,r21_89,r21_90,r21_91,r21_92,r21_93,r21_94,r21_95,r21_96,
		r21_97,r21_98,r21_99,r21_100,r21_101,r21_102,r21_103,r21_104,r21_105,r21_106,r21_107,r21_108,r21_109,r21_110,r21_111,r21_112,
		r21_113,r21_114,r21_115,r21_116,r21_117,r21_118,r21_119,r21_120,r21_121,r21_122,r21_123,r21_124,r21_125,r21_126,
	r22_0,r22_1,r22_2,r22_3,r22_4,r22_5,r22_6,r22_7,r22_8,r22_9,r22_10,r22_11,r22_12,r22_13,r22_14,r22_15,r22_16,
		r22_17,r22_18,r22_19,r22_20,r22_21,r22_22,r22_23,r22_24,r22_25,r22_26,r22_27,r22_28,r22_29,r22_30,r22_31,r22_32,
		r22_33,r22_34,r22_35,r22_36,r22_37,r22_38,r22_39,r22_40,r22_41,r22_42,r22_43,r22_44,r22_45,r22_46,r22_47,r22_48,
		r22_49,r22_50,r22_51,r22_52,r22_53,r22_54,r22_55,r22_56,r22_57,r22_58,r22_59,r22_60,r22_61,r22_62,r22_63,r22_64,
		r22_65,r22_66,r22_67,r22_68,r22_69,r22_70,r22_71,r22_72,r22_73,r22_74,r22_75,r22_76,r22_77,r22_78,r22_79,r22_80,
		r22_81,r22_82,r22_83,r22_84,r22_85,r22_86,r22_87,r22_88,r22_89,r22_90,r22_91,r22_92,r22_93,r22_94,r22_95,r22_96,
		r22_97,r22_98,r22_99,r22_100,r22_101,r22_102,r22_103,r22_104,r22_105,r22_106,r22_107,r22_108,r22_109,r22_110,r22_111,r22_112,
		r22_113,r22_114,r22_115,r22_116,r22_117,r22_118,r22_119,r22_120,r22_121,r22_122,r22_123,r22_124,r22_125,r22_126,
	r23_0,r23_1,r23_2,r23_3,r23_4,r23_5,r23_6,r23_7,r23_8,r23_9,r23_10,r23_11,r23_12,r23_13,r23_14,r23_15,r23_16,
		r23_17,r23_18,r23_19,r23_20,r23_21,r23_22,r23_23,r23_24,r23_25,r23_26,r23_27,r23_28,r23_29,r23_30,r23_31,r23_32,
		r23_33,r23_34,r23_35,r23_36,r23_37,r23_38,r23_39,r23_40,r23_41,r23_42,r23_43,r23_44,r23_45,r23_46,r23_47,r23_48,
		r23_49,r23_50,r23_51,r23_52,r23_53,r23_54,r23_55,r23_56,r23_57,r23_58,r23_59,r23_60,r23_61,r23_62,r23_63,r23_64,
		r23_65,r23_66,r23_67,r23_68,r23_69,r23_70,r23_71,r23_72,r23_73,r23_74,r23_75,r23_76,r23_77,r23_78,r23_79,r23_80,
		r23_81,r23_82,r23_83,r23_84,r23_85,r23_86,r23_87,r23_88,r23_89,r23_90,r23_91,r23_92,r23_93,r23_94,r23_95,r23_96,
		r23_97,r23_98,r23_99,r23_100,r23_101,r23_102,r23_103,r23_104,r23_105,r23_106,r23_107,r23_108,r23_109,r23_110,r23_111,r23_112,
		r23_113,r23_114,r23_115,r23_116,r23_117,r23_118,r23_119,r23_120,r23_121,r23_122,r23_123,r23_124,r23_125,r23_126,
	r24_0,r24_1,r24_2,r24_3,r24_4,r24_5,r24_6,r24_7,r24_8,r24_9,r24_10,r24_11,r24_12,r24_13,r24_14,r24_15,r24_16,
		r24_17,r24_18,r24_19,r24_20,r24_21,r24_22,r24_23,r24_24,r24_25,r24_26,r24_27,r24_28,r24_29,r24_30,r24_31,r24_32,
		r24_33,r24_34,r24_35,r24_36,r24_37,r24_38,r24_39,r24_40,r24_41,r24_42,r24_43,r24_44,r24_45,r24_46,r24_47,r24_48,
		r24_49,r24_50,r24_51,r24_52,r24_53,r24_54,r24_55,r24_56,r24_57,r24_58,r24_59,r24_60,r24_61,r24_62,r24_63,r24_64,
		r24_65,r24_66,r24_67,r24_68,r24_69,r24_70,r24_71,r24_72,r24_73,r24_74,r24_75,r24_76,r24_77,r24_78,r24_79,r24_80,
		r24_81,r24_82,r24_83,r24_84,r24_85,r24_86,r24_87,r24_88,r24_89,r24_90,r24_91,r24_92,r24_93,r24_94,r24_95,r24_96,
		r24_97,r24_98,r24_99,r24_100,r24_101,r24_102,r24_103,r24_104,r24_105,r24_106,r24_107,r24_108,r24_109,r24_110,r24_111,r24_112,
		r24_113,r24_114,r24_115,r24_116,r24_117,r24_118,r24_119,r24_120,r24_121,r24_122,r24_123,r24_124,r24_125,r24_126,
	r25_0,r25_1,r25_2,r25_3,r25_4,r25_5,r25_6,r25_7,r25_8,r25_9,r25_10,r25_11,r25_12,r25_13,r25_14,r25_15,r25_16,
		r25_17,r25_18,r25_19,r25_20,r25_21,r25_22,r25_23,r25_24,r25_25,r25_26,r25_27,r25_28,r25_29,r25_30,r25_31,r25_32,
		r25_33,r25_34,r25_35,r25_36,r25_37,r25_38,r25_39,r25_40,r25_41,r25_42,r25_43,r25_44,r25_45,r25_46,r25_47,r25_48,
		r25_49,r25_50,r25_51,r25_52,r25_53,r25_54,r25_55,r25_56,r25_57,r25_58,r25_59,r25_60,r25_61,r25_62,r25_63,r25_64,
		r25_65,r25_66,r25_67,r25_68,r25_69,r25_70,r25_71,r25_72,r25_73,r25_74,r25_75,r25_76,r25_77,r25_78,r25_79,r25_80,
		r25_81,r25_82,r25_83,r25_84,r25_85,r25_86,r25_87,r25_88,r25_89,r25_90,r25_91,r25_92,r25_93,r25_94,r25_95,r25_96,
		r25_97,r25_98,r25_99,r25_100,r25_101,r25_102,r25_103,r25_104,r25_105,r25_106,r25_107,r25_108,r25_109,r25_110,r25_111,r25_112,
		r25_113,r25_114,r25_115,r25_116,r25_117,r25_118,r25_119,r25_120,r25_121,r25_122,r25_123,r25_124,r25_125,r25_126,
	r26_0,r26_1,r26_2,r26_3,r26_4,r26_5,r26_6,r26_7,r26_8,r26_9,r26_10,r26_11,r26_12,r26_13,r26_14,r26_15,r26_16,
		r26_17,r26_18,r26_19,r26_20,r26_21,r26_22,r26_23,r26_24,r26_25,r26_26,r26_27,r26_28,r26_29,r26_30,r26_31,r26_32,
		r26_33,r26_34,r26_35,r26_36,r26_37,r26_38,r26_39,r26_40,r26_41,r26_42,r26_43,r26_44,r26_45,r26_46,r26_47,r26_48,
		r26_49,r26_50,r26_51,r26_52,r26_53,r26_54,r26_55,r26_56,r26_57,r26_58,r26_59,r26_60,r26_61,r26_62,r26_63,r26_64,
		r26_65,r26_66,r26_67,r26_68,r26_69,r26_70,r26_71,r26_72,r26_73,r26_74,r26_75,r26_76,r26_77,r26_78,r26_79,r26_80,
		r26_81,r26_82,r26_83,r26_84,r26_85,r26_86,r26_87,r26_88,r26_89,r26_90,r26_91,r26_92,r26_93,r26_94,r26_95,r26_96,
		r26_97,r26_98,r26_99,r26_100,r26_101,r26_102,r26_103,r26_104,r26_105,r26_106,r26_107,r26_108,r26_109,r26_110,r26_111,r26_112,
		r26_113,r26_114,r26_115,r26_116,r26_117,r26_118,r26_119,r26_120,r26_121,r26_122,r26_123,r26_124,r26_125,r26_126,
	r27_0,r27_1,r27_2,r27_3,r27_4,r27_5,r27_6,r27_7,r27_8,r27_9,r27_10,r27_11,r27_12,r27_13,r27_14,r27_15,r27_16,
		r27_17,r27_18,r27_19,r27_20,r27_21,r27_22,r27_23,r27_24,r27_25,r27_26,r27_27,r27_28,r27_29,r27_30,r27_31,r27_32,
		r27_33,r27_34,r27_35,r27_36,r27_37,r27_38,r27_39,r27_40,r27_41,r27_42,r27_43,r27_44,r27_45,r27_46,r27_47,r27_48,
		r27_49,r27_50,r27_51,r27_52,r27_53,r27_54,r27_55,r27_56,r27_57,r27_58,r27_59,r27_60,r27_61,r27_62,r27_63,r27_64,
		r27_65,r27_66,r27_67,r27_68,r27_69,r27_70,r27_71,r27_72,r27_73,r27_74,r27_75,r27_76,r27_77,r27_78,r27_79,r27_80,
		r27_81,r27_82,r27_83,r27_84,r27_85,r27_86,r27_87,r27_88,r27_89,r27_90,r27_91,r27_92,r27_93,r27_94,r27_95,r27_96,
		r27_97,r27_98,r27_99,r27_100,r27_101,r27_102,r27_103,r27_104,r27_105,r27_106,r27_107,r27_108,r27_109,r27_110,r27_111,r27_112,
		r27_113,r27_114,r27_115,r27_116,r27_117,r27_118,r27_119,r27_120,r27_121,r27_122,r27_123,r27_124,r27_125,r27_126,
	r28_0,r28_1,r28_2,r28_3,r28_4,r28_5,r28_6,r28_7,r28_8,r28_9,r28_10,r28_11,r28_12,r28_13,r28_14,r28_15,r28_16,
		r28_17,r28_18,r28_19,r28_20,r28_21,r28_22,r28_23,r28_24,r28_25,r28_26,r28_27,r28_28,r28_29,r28_30,r28_31,r28_32,
		r28_33,r28_34,r28_35,r28_36,r28_37,r28_38,r28_39,r28_40,r28_41,r28_42,r28_43,r28_44,r28_45,r28_46,r28_47,r28_48,
		r28_49,r28_50,r28_51,r28_52,r28_53,r28_54,r28_55,r28_56,r28_57,r28_58,r28_59,r28_60,r28_61,r28_62,r28_63,r28_64,
		r28_65,r28_66,r28_67,r28_68,r28_69,r28_70,r28_71,r28_72,r28_73,r28_74,r28_75,r28_76,r28_77,r28_78,r28_79,r28_80,
		r28_81,r28_82,r28_83,r28_84,r28_85,r28_86,r28_87,r28_88,r28_89,r28_90,r28_91,r28_92,r28_93,r28_94,r28_95,r28_96,
		r28_97,r28_98,r28_99,r28_100,r28_101,r28_102,r28_103,r28_104,r28_105,r28_106,r28_107,r28_108,r28_109,r28_110,r28_111,r28_112,
		r28_113,r28_114,r28_115,r28_116,r28_117,r28_118,r28_119,r28_120,r28_121,r28_122,r28_123,r28_124,r28_125,r28_126,
	r29_0,r29_1,r29_2,r29_3,r29_4,r29_5,r29_6,r29_7,r29_8,r29_9,r29_10,r29_11,r29_12,r29_13,r29_14,r29_15,r29_16,
		r29_17,r29_18,r29_19,r29_20,r29_21,r29_22,r29_23,r29_24,r29_25,r29_26,r29_27,r29_28,r29_29,r29_30,r29_31,r29_32,
		r29_33,r29_34,r29_35,r29_36,r29_37,r29_38,r29_39,r29_40,r29_41,r29_42,r29_43,r29_44,r29_45,r29_46,r29_47,r29_48,
		r29_49,r29_50,r29_51,r29_52,r29_53,r29_54,r29_55,r29_56,r29_57,r29_58,r29_59,r29_60,r29_61,r29_62,r29_63,r29_64,
		r29_65,r29_66,r29_67,r29_68,r29_69,r29_70,r29_71,r29_72,r29_73,r29_74,r29_75,r29_76,r29_77,r29_78,r29_79,r29_80,
		r29_81,r29_82,r29_83,r29_84,r29_85,r29_86,r29_87,r29_88,r29_89,r29_90,r29_91,r29_92,r29_93,r29_94,r29_95,r29_96,
		r29_97,r29_98,r29_99,r29_100,r29_101,r29_102,r29_103,r29_104,r29_105,r29_106,r29_107,r29_108,r29_109,r29_110,r29_111,r29_112,
		r29_113,r29_114,r29_115,r29_116,r29_117,r29_118,r29_119,r29_120,r29_121,r29_122,r29_123,r29_124,r29_125,r29_126,
	r30_0,r30_1,r30_2,r30_3,r30_4,r30_5,r30_6,r30_7,r30_8,r30_9,r30_10,r30_11,r30_12,r30_13,r30_14,r30_15,r30_16,
		r30_17,r30_18,r30_19,r30_20,r30_21,r30_22,r30_23,r30_24,r30_25,r30_26,r30_27,r30_28,r30_29,r30_30,r30_31,r30_32,
		r30_33,r30_34,r30_35,r30_36,r30_37,r30_38,r30_39,r30_40,r30_41,r30_42,r30_43,r30_44,r30_45,r30_46,r30_47,r30_48,
		r30_49,r30_50,r30_51,r30_52,r30_53,r30_54,r30_55,r30_56,r30_57,r30_58,r30_59,r30_60,r30_61,r30_62,r30_63,r30_64,
		r30_65,r30_66,r30_67,r30_68,r30_69,r30_70,r30_71,r30_72,r30_73,r30_74,r30_75,r30_76,r30_77,r30_78,r30_79,r30_80,
		r30_81,r30_82,r30_83,r30_84,r30_85,r30_86,r30_87,r30_88,r30_89,r30_90,r30_91,r30_92,r30_93,r30_94,r30_95,r30_96,
		r30_97,r30_98,r30_99,r30_100,r30_101,r30_102,r30_103,r30_104,r30_105,r30_106,r30_107,r30_108,r30_109,r30_110,r30_111,r30_112,
		r30_113,r30_114,r30_115,r30_116,r30_117,r30_118,r30_119,r30_120,r30_121,r30_122,r30_123,r30_124,r30_125,r30_126,
	r31_0,r31_1,r31_2,r31_3,r31_4,r31_5,r31_6,r31_7,r31_8,r31_9,r31_10,r31_11,r31_12,r31_13,r31_14,r31_15,r31_16,
		r31_17,r31_18,r31_19,r31_20,r31_21,r31_22,r31_23,r31_24,r31_25,r31_26,r31_27,r31_28,r31_29,r31_30,r31_31,r31_32,
		r31_33,r31_34,r31_35,r31_36,r31_37,r31_38,r31_39,r31_40,r31_41,r31_42,r31_43,r31_44,r31_45,r31_46,r31_47,r31_48,
		r31_49,r31_50,r31_51,r31_52,r31_53,r31_54,r31_55,r31_56,r31_57,r31_58,r31_59,r31_60,r31_61,r31_62,r31_63,r31_64,
		r31_65,r31_66,r31_67,r31_68,r31_69,r31_70,r31_71,r31_72,r31_73,r31_74,r31_75,r31_76,r31_77,r31_78,r31_79,r31_80,
		r31_81,r31_82,r31_83,r31_84,r31_85,r31_86,r31_87,r31_88,r31_89,r31_90,r31_91,r31_92,r31_93,r31_94,r31_95,r31_96,
		r31_97,r31_98,r31_99,r31_100,r31_101,r31_102,r31_103,r31_104,r31_105,r31_106,r31_107,r31_108,r31_109,r31_110,r31_111,r31_112,
		r31_113,r31_114,r31_115,r31_116,r31_117,r31_118,r31_119,r31_120,r31_121,r31_122,r31_123,r31_124,r31_125,r31_126,
	r32_0,r32_1,r32_2,r32_3,r32_4,r32_5,r32_6,r32_7,r32_8,r32_9,r32_10,r32_11,r32_12,r32_13,r32_14,r32_15,r32_16,
		r32_17,r32_18,r32_19,r32_20,r32_21,r32_22,r32_23,r32_24,r32_25,r32_26,r32_27,r32_28,r32_29,r32_30,r32_31,r32_32,
		r32_33,r32_34,r32_35,r32_36,r32_37,r32_38,r32_39,r32_40,r32_41,r32_42,r32_43,r32_44,r32_45,r32_46,r32_47,r32_48,
		r32_49,r32_50,r32_51,r32_52,r32_53,r32_54,r32_55,r32_56,r32_57,r32_58,r32_59,r32_60,r32_61,r32_62,r32_63,r32_64,
		r32_65,r32_66,r32_67,r32_68,r32_69,r32_70,r32_71,r32_72,r32_73,r32_74,r32_75,r32_76,r32_77,r32_78,r32_79,r32_80,
		r32_81,r32_82,r32_83,r32_84,r32_85,r32_86,r32_87,r32_88,r32_89,r32_90,r32_91,r32_92,r32_93,r32_94,r32_95,r32_96,
		r32_97,r32_98,r32_99,r32_100,r32_101,r32_102,r32_103,r32_104,r32_105,r32_106,r32_107,r32_108,r32_109,r32_110,r32_111,r32_112,
		r32_113,r32_114,r32_115,r32_116,r32_117,r32_118,r32_119,r32_120,r32_121,r32_122,r32_123,r32_124,r32_125,r32_126,
	r33_0,r33_1,r33_2,r33_3,r33_4,r33_5,r33_6,r33_7,r33_8,r33_9,r33_10,r33_11,r33_12,r33_13,r33_14,r33_15,r33_16,
		r33_17,r33_18,r33_19,r33_20,r33_21,r33_22,r33_23,r33_24,r33_25,r33_26,r33_27,r33_28,r33_29,r33_30,r33_31,r33_32,
		r33_33,r33_34,r33_35,r33_36,r33_37,r33_38,r33_39,r33_40,r33_41,r33_42,r33_43,r33_44,r33_45,r33_46,r33_47,r33_48,
		r33_49,r33_50,r33_51,r33_52,r33_53,r33_54,r33_55,r33_56,r33_57,r33_58,r33_59,r33_60,r33_61,r33_62,r33_63,r33_64,
		r33_65,r33_66,r33_67,r33_68,r33_69,r33_70,r33_71,r33_72,r33_73,r33_74,r33_75,r33_76,r33_77,r33_78,r33_79,r33_80,
		r33_81,r33_82,r33_83,r33_84,r33_85,r33_86,r33_87,r33_88,r33_89,r33_90,r33_91,r33_92,r33_93,r33_94,r33_95,r33_96,
		r33_97,r33_98,r33_99,r33_100,r33_101,r33_102,r33_103,r33_104,r33_105,r33_106,r33_107,r33_108,r33_109,r33_110,r33_111,r33_112,
		r33_113,r33_114,r33_115,r33_116,r33_117,r33_118,r33_119,r33_120,r33_121,r33_122,r33_123,r33_124,r33_125,r33_126,
	r34_0,r34_1,r34_2,r34_3,r34_4,r34_5,r34_6,r34_7,r34_8,r34_9,r34_10,r34_11,r34_12,r34_13,r34_14,r34_15,r34_16,
		r34_17,r34_18,r34_19,r34_20,r34_21,r34_22,r34_23,r34_24,r34_25,r34_26,r34_27,r34_28,r34_29,r34_30,r34_31,r34_32,
		r34_33,r34_34,r34_35,r34_36,r34_37,r34_38,r34_39,r34_40,r34_41,r34_42,r34_43,r34_44,r34_45,r34_46,r34_47,r34_48,
		r34_49,r34_50,r34_51,r34_52,r34_53,r34_54,r34_55,r34_56,r34_57,r34_58,r34_59,r34_60,r34_61,r34_62,r34_63,r34_64,
		r34_65,r34_66,r34_67,r34_68,r34_69,r34_70,r34_71,r34_72,r34_73,r34_74,r34_75,r34_76,r34_77,r34_78,r34_79,r34_80,
		r34_81,r34_82,r34_83,r34_84,r34_85,r34_86,r34_87,r34_88,r34_89,r34_90,r34_91,r34_92,r34_93,r34_94,r34_95,r34_96,
		r34_97,r34_98,r34_99,r34_100,r34_101,r34_102,r34_103,r34_104,r34_105,r34_106,r34_107,r34_108,r34_109,r34_110,r34_111,r34_112,
		r34_113,r34_114,r34_115,r34_116,r34_117,r34_118,r34_119,r34_120,r34_121,r34_122,r34_123,r34_124,r34_125,r34_126,
	r35_0,r35_1,r35_2,r35_3,r35_4,r35_5,r35_6,r35_7,r35_8,r35_9,r35_10,r35_11,r35_12,r35_13,r35_14,r35_15,r35_16,
		r35_17,r35_18,r35_19,r35_20,r35_21,r35_22,r35_23,r35_24,r35_25,r35_26,r35_27,r35_28,r35_29,r35_30,r35_31,r35_32,
		r35_33,r35_34,r35_35,r35_36,r35_37,r35_38,r35_39,r35_40,r35_41,r35_42,r35_43,r35_44,r35_45,r35_46,r35_47,r35_48,
		r35_49,r35_50,r35_51,r35_52,r35_53,r35_54,r35_55,r35_56,r35_57,r35_58,r35_59,r35_60,r35_61,r35_62,r35_63,r35_64,
		r35_65,r35_66,r35_67,r35_68,r35_69,r35_70,r35_71,r35_72,r35_73,r35_74,r35_75,r35_76,r35_77,r35_78,r35_79,r35_80,
		r35_81,r35_82,r35_83,r35_84,r35_85,r35_86,r35_87,r35_88,r35_89,r35_90,r35_91,r35_92,r35_93,r35_94,r35_95,r35_96,
		r35_97,r35_98,r35_99,r35_100,r35_101,r35_102,r35_103,r35_104,r35_105,r35_106,r35_107,r35_108,r35_109,r35_110,r35_111,r35_112,
		r35_113,r35_114,r35_115,r35_116,r35_117,r35_118,r35_119,r35_120,r35_121,r35_122,r35_123,r35_124,r35_125,r35_126,
	r36_0,r36_1,r36_2,r36_3,r36_4,r36_5,r36_6,r36_7,r36_8,r36_9,r36_10,r36_11,r36_12,r36_13,r36_14,r36_15,r36_16,
		r36_17,r36_18,r36_19,r36_20,r36_21,r36_22,r36_23,r36_24,r36_25,r36_26,r36_27,r36_28,r36_29,r36_30,r36_31,r36_32,
		r36_33,r36_34,r36_35,r36_36,r36_37,r36_38,r36_39,r36_40,r36_41,r36_42,r36_43,r36_44,r36_45,r36_46,r36_47,r36_48,
		r36_49,r36_50,r36_51,r36_52,r36_53,r36_54,r36_55,r36_56,r36_57,r36_58,r36_59,r36_60,r36_61,r36_62,r36_63,r36_64,
		r36_65,r36_66,r36_67,r36_68,r36_69,r36_70,r36_71,r36_72,r36_73,r36_74,r36_75,r36_76,r36_77,r36_78,r36_79,r36_80,
		r36_81,r36_82,r36_83,r36_84,r36_85,r36_86,r36_87,r36_88,r36_89,r36_90,r36_91,r36_92,r36_93,r36_94,r36_95,r36_96,
		r36_97,r36_98,r36_99,r36_100,r36_101,r36_102,r36_103,r36_104,r36_105,r36_106,r36_107,r36_108,r36_109,r36_110,r36_111,r36_112,
		r36_113,r36_114,r36_115,r36_116,r36_117,r36_118,r36_119,r36_120,r36_121,r36_122,r36_123,r36_124,r36_125,r36_126,
	r37_0,r37_1,r37_2,r37_3,r37_4,r37_5,r37_6,r37_7,r37_8,r37_9,r37_10,r37_11,r37_12,r37_13,r37_14,r37_15,r37_16,
		r37_17,r37_18,r37_19,r37_20,r37_21,r37_22,r37_23,r37_24,r37_25,r37_26,r37_27,r37_28,r37_29,r37_30,r37_31,r37_32,
		r37_33,r37_34,r37_35,r37_36,r37_37,r37_38,r37_39,r37_40,r37_41,r37_42,r37_43,r37_44,r37_45,r37_46,r37_47,r37_48,
		r37_49,r37_50,r37_51,r37_52,r37_53,r37_54,r37_55,r37_56,r37_57,r37_58,r37_59,r37_60,r37_61,r37_62,r37_63,r37_64,
		r37_65,r37_66,r37_67,r37_68,r37_69,r37_70,r37_71,r37_72,r37_73,r37_74,r37_75,r37_76,r37_77,r37_78,r37_79,r37_80,
		r37_81,r37_82,r37_83,r37_84,r37_85,r37_86,r37_87,r37_88,r37_89,r37_90,r37_91,r37_92,r37_93,r37_94,r37_95,r37_96,
		r37_97,r37_98,r37_99,r37_100,r37_101,r37_102,r37_103,r37_104,r37_105,r37_106,r37_107,r37_108,r37_109,r37_110,r37_111,r37_112,
		r37_113,r37_114,r37_115,r37_116,r37_117,r37_118,r37_119,r37_120,r37_121,r37_122,r37_123,r37_124,r37_125,r37_126,
	r38_0,r38_1,r38_2,r38_3,r38_4,r38_5,r38_6,r38_7,r38_8,r38_9,r38_10,r38_11,r38_12,r38_13,r38_14,r38_15,r38_16,
		r38_17,r38_18,r38_19,r38_20,r38_21,r38_22,r38_23,r38_24,r38_25,r38_26,r38_27,r38_28,r38_29,r38_30,r38_31,r38_32,
		r38_33,r38_34,r38_35,r38_36,r38_37,r38_38,r38_39,r38_40,r38_41,r38_42,r38_43,r38_44,r38_45,r38_46,r38_47,r38_48,
		r38_49,r38_50,r38_51,r38_52,r38_53,r38_54,r38_55,r38_56,r38_57,r38_58,r38_59,r38_60,r38_61,r38_62,r38_63,r38_64,
		r38_65,r38_66,r38_67,r38_68,r38_69,r38_70,r38_71,r38_72,r38_73,r38_74,r38_75,r38_76,r38_77,r38_78,r38_79,r38_80,
		r38_81,r38_82,r38_83,r38_84,r38_85,r38_86,r38_87,r38_88,r38_89,r38_90,r38_91,r38_92,r38_93,r38_94,r38_95,r38_96,
		r38_97,r38_98,r38_99,r38_100,r38_101,r38_102,r38_103,r38_104,r38_105,r38_106,r38_107,r38_108,r38_109,r38_110,r38_111,r38_112,
		r38_113,r38_114,r38_115,r38_116,r38_117,r38_118,r38_119,r38_120,r38_121,r38_122,r38_123,r38_124,r38_125,r38_126,
	r39_0,r39_1,r39_2,r39_3,r39_4,r39_5,r39_6,r39_7,r39_8,r39_9,r39_10,r39_11,r39_12,r39_13,r39_14,r39_15,r39_16,
		r39_17,r39_18,r39_19,r39_20,r39_21,r39_22,r39_23,r39_24,r39_25,r39_26,r39_27,r39_28,r39_29,r39_30,r39_31,r39_32,
		r39_33,r39_34,r39_35,r39_36,r39_37,r39_38,r39_39,r39_40,r39_41,r39_42,r39_43,r39_44,r39_45,r39_46,r39_47,r39_48,
		r39_49,r39_50,r39_51,r39_52,r39_53,r39_54,r39_55,r39_56,r39_57,r39_58,r39_59,r39_60,r39_61,r39_62,r39_63,r39_64,
		r39_65,r39_66,r39_67,r39_68,r39_69,r39_70,r39_71,r39_72,r39_73,r39_74,r39_75,r39_76,r39_77,r39_78,r39_79,r39_80,
		r39_81,r39_82,r39_83,r39_84,r39_85,r39_86,r39_87,r39_88,r39_89,r39_90,r39_91,r39_92,r39_93,r39_94,r39_95,r39_96,
		r39_97,r39_98,r39_99,r39_100,r39_101,r39_102,r39_103,r39_104,r39_105,r39_106,r39_107,r39_108,r39_109,r39_110,r39_111,r39_112,
		r39_113,r39_114,r39_115,r39_116,r39_117,r39_118,r39_119,r39_120,r39_121,r39_122,r39_123,r39_124,r39_125,r39_126,
	r40_0,r40_1,r40_2,r40_3,r40_4,r40_5,r40_6,r40_7,r40_8,r40_9,r40_10,r40_11,r40_12,r40_13,r40_14,r40_15,r40_16,
		r40_17,r40_18,r40_19,r40_20,r40_21,r40_22,r40_23,r40_24,r40_25,r40_26,r40_27,r40_28,r40_29,r40_30,r40_31,r40_32,
		r40_33,r40_34,r40_35,r40_36,r40_37,r40_38,r40_39,r40_40,r40_41,r40_42,r40_43,r40_44,r40_45,r40_46,r40_47,r40_48,
		r40_49,r40_50,r40_51,r40_52,r40_53,r40_54,r40_55,r40_56,r40_57,r40_58,r40_59,r40_60,r40_61,r40_62,r40_63,r40_64,
		r40_65,r40_66,r40_67,r40_68,r40_69,r40_70,r40_71,r40_72,r40_73,r40_74,r40_75,r40_76,r40_77,r40_78,r40_79,r40_80,
		r40_81,r40_82,r40_83,r40_84,r40_85,r40_86,r40_87,r40_88,r40_89,r40_90,r40_91,r40_92,r40_93,r40_94,r40_95,r40_96,
		r40_97,r40_98,r40_99,r40_100,r40_101,r40_102,r40_103,r40_104,r40_105,r40_106,r40_107,r40_108,r40_109,r40_110,r40_111,r40_112,
		r40_113,r40_114,r40_115,r40_116,r40_117,r40_118,r40_119,r40_120,r40_121,r40_122,r40_123,r40_124,r40_125,r40_126,
	r41_0,r41_1,r41_2,r41_3,r41_4,r41_5,r41_6,r41_7,r41_8,r41_9,r41_10,r41_11,r41_12,r41_13,r41_14,r41_15,r41_16,
		r41_17,r41_18,r41_19,r41_20,r41_21,r41_22,r41_23,r41_24,r41_25,r41_26,r41_27,r41_28,r41_29,r41_30,r41_31,r41_32,
		r41_33,r41_34,r41_35,r41_36,r41_37,r41_38,r41_39,r41_40,r41_41,r41_42,r41_43,r41_44,r41_45,r41_46,r41_47,r41_48,
		r41_49,r41_50,r41_51,r41_52,r41_53,r41_54,r41_55,r41_56,r41_57,r41_58,r41_59,r41_60,r41_61,r41_62,r41_63,r41_64,
		r41_65,r41_66,r41_67,r41_68,r41_69,r41_70,r41_71,r41_72,r41_73,r41_74,r41_75,r41_76,r41_77,r41_78,r41_79,r41_80,
		r41_81,r41_82,r41_83,r41_84,r41_85,r41_86,r41_87,r41_88,r41_89,r41_90,r41_91,r41_92,r41_93,r41_94,r41_95,r41_96,
		r41_97,r41_98,r41_99,r41_100,r41_101,r41_102,r41_103,r41_104,r41_105,r41_106,r41_107,r41_108,r41_109,r41_110,r41_111,r41_112,
		r41_113,r41_114,r41_115,r41_116,r41_117,r41_118,r41_119,r41_120,r41_121,r41_122,r41_123,r41_124,r41_125,r41_126,
	r42_0,r42_1,r42_2,r42_3,r42_4,r42_5,r42_6,r42_7,r42_8,r42_9,r42_10,r42_11,r42_12,r42_13,r42_14,r42_15,r42_16,
		r42_17,r42_18,r42_19,r42_20,r42_21,r42_22,r42_23,r42_24,r42_25,r42_26,r42_27,r42_28,r42_29,r42_30,r42_31,r42_32,
		r42_33,r42_34,r42_35,r42_36,r42_37,r42_38,r42_39,r42_40,r42_41,r42_42,r42_43,r42_44,r42_45,r42_46,r42_47,r42_48,
		r42_49,r42_50,r42_51,r42_52,r42_53,r42_54,r42_55,r42_56,r42_57,r42_58,r42_59,r42_60,r42_61,r42_62,r42_63,r42_64,
		r42_65,r42_66,r42_67,r42_68,r42_69,r42_70,r42_71,r42_72,r42_73,r42_74,r42_75,r42_76,r42_77,r42_78,r42_79,r42_80,
		r42_81,r42_82,r42_83,r42_84,r42_85,r42_86,r42_87,r42_88,r42_89,r42_90,r42_91,r42_92,r42_93,r42_94,r42_95,r42_96,
		r42_97,r42_98,r42_99,r42_100,r42_101,r42_102,r42_103,r42_104,r42_105,r42_106,r42_107,r42_108,r42_109,r42_110,r42_111,r42_112,
		r42_113,r42_114,r42_115,r42_116,r42_117,r42_118,r42_119,r42_120,r42_121,r42_122,r42_123,r42_124,r42_125,r42_126,
	r43_0,r43_1,r43_2,r43_3,r43_4,r43_5,r43_6,r43_7,r43_8,r43_9,r43_10,r43_11,r43_12,r43_13,r43_14,r43_15,r43_16,
		r43_17,r43_18,r43_19,r43_20,r43_21,r43_22,r43_23,r43_24,r43_25,r43_26,r43_27,r43_28,r43_29,r43_30,r43_31,r43_32,
		r43_33,r43_34,r43_35,r43_36,r43_37,r43_38,r43_39,r43_40,r43_41,r43_42,r43_43,r43_44,r43_45,r43_46,r43_47,r43_48,
		r43_49,r43_50,r43_51,r43_52,r43_53,r43_54,r43_55,r43_56,r43_57,r43_58,r43_59,r43_60,r43_61,r43_62,r43_63,r43_64,
		r43_65,r43_66,r43_67,r43_68,r43_69,r43_70,r43_71,r43_72,r43_73,r43_74,r43_75,r43_76,r43_77,r43_78,r43_79,r43_80,
		r43_81,r43_82,r43_83,r43_84,r43_85,r43_86,r43_87,r43_88,r43_89,r43_90,r43_91,r43_92,r43_93,r43_94,r43_95,r43_96,
		r43_97,r43_98,r43_99,r43_100,r43_101,r43_102,r43_103,r43_104,r43_105,r43_106,r43_107,r43_108,r43_109,r43_110,r43_111,r43_112,
		r43_113,r43_114,r43_115,r43_116,r43_117,r43_118,r43_119,r43_120,r43_121,r43_122,r43_123,r43_124,r43_125,r43_126,
	r44_0,r44_1,r44_2,r44_3,r44_4,r44_5,r44_6,r44_7,r44_8,r44_9,r44_10,r44_11,r44_12,r44_13,r44_14,r44_15,r44_16,
		r44_17,r44_18,r44_19,r44_20,r44_21,r44_22,r44_23,r44_24,r44_25,r44_26,r44_27,r44_28,r44_29,r44_30,r44_31,r44_32,
		r44_33,r44_34,r44_35,r44_36,r44_37,r44_38,r44_39,r44_40,r44_41,r44_42,r44_43,r44_44,r44_45,r44_46,r44_47,r44_48,
		r44_49,r44_50,r44_51,r44_52,r44_53,r44_54,r44_55,r44_56,r44_57,r44_58,r44_59,r44_60,r44_61,r44_62,r44_63,r44_64,
		r44_65,r44_66,r44_67,r44_68,r44_69,r44_70,r44_71,r44_72,r44_73,r44_74,r44_75,r44_76,r44_77,r44_78,r44_79,r44_80,
		r44_81,r44_82,r44_83,r44_84,r44_85,r44_86,r44_87,r44_88,r44_89,r44_90,r44_91,r44_92,r44_93,r44_94,r44_95,r44_96,
		r44_97,r44_98,r44_99,r44_100,r44_101,r44_102,r44_103,r44_104,r44_105,r44_106,r44_107,r44_108,r44_109,r44_110,r44_111,r44_112,
		r44_113,r44_114,r44_115,r44_116,r44_117,r44_118,r44_119,r44_120,r44_121,r44_122,r44_123,r44_124,r44_125,r44_126,
	r45_0,r45_1,r45_2,r45_3,r45_4,r45_5,r45_6,r45_7,r45_8,r45_9,r45_10,r45_11,r45_12,r45_13,r45_14,r45_15,r45_16,
		r45_17,r45_18,r45_19,r45_20,r45_21,r45_22,r45_23,r45_24,r45_25,r45_26,r45_27,r45_28,r45_29,r45_30,r45_31,r45_32,
		r45_33,r45_34,r45_35,r45_36,r45_37,r45_38,r45_39,r45_40,r45_41,r45_42,r45_43,r45_44,r45_45,r45_46,r45_47,r45_48,
		r45_49,r45_50,r45_51,r45_52,r45_53,r45_54,r45_55,r45_56,r45_57,r45_58,r45_59,r45_60,r45_61,r45_62,r45_63,r45_64,
		r45_65,r45_66,r45_67,r45_68,r45_69,r45_70,r45_71,r45_72,r45_73,r45_74,r45_75,r45_76,r45_77,r45_78,r45_79,r45_80,
		r45_81,r45_82,r45_83,r45_84,r45_85,r45_86,r45_87,r45_88,r45_89,r45_90,r45_91,r45_92,r45_93,r45_94,r45_95,r45_96,
		r45_97,r45_98,r45_99,r45_100,r45_101,r45_102,r45_103,r45_104,r45_105,r45_106,r45_107,r45_108,r45_109,r45_110,r45_111,r45_112,
		r45_113,r45_114,r45_115,r45_116,r45_117,r45_118,r45_119,r45_120,r45_121,r45_122,r45_123,r45_124,r45_125,r45_126,
	r46_0,r46_1,r46_2,r46_3,r46_4,r46_5,r46_6,r46_7,r46_8,r46_9,r46_10,r46_11,r46_12,r46_13,r46_14,r46_15,r46_16,
		r46_17,r46_18,r46_19,r46_20,r46_21,r46_22,r46_23,r46_24,r46_25,r46_26,r46_27,r46_28,r46_29,r46_30,r46_31,r46_32,
		r46_33,r46_34,r46_35,r46_36,r46_37,r46_38,r46_39,r46_40,r46_41,r46_42,r46_43,r46_44,r46_45,r46_46,r46_47,r46_48,
		r46_49,r46_50,r46_51,r46_52,r46_53,r46_54,r46_55,r46_56,r46_57,r46_58,r46_59,r46_60,r46_61,r46_62,r46_63,r46_64,
		r46_65,r46_66,r46_67,r46_68,r46_69,r46_70,r46_71,r46_72,r46_73,r46_74,r46_75,r46_76,r46_77,r46_78,r46_79,r46_80,
		r46_81,r46_82,r46_83,r46_84,r46_85,r46_86,r46_87,r46_88,r46_89,r46_90,r46_91,r46_92,r46_93,r46_94,r46_95,r46_96,
		r46_97,r46_98,r46_99,r46_100,r46_101,r46_102,r46_103,r46_104,r46_105,r46_106,r46_107,r46_108,r46_109,r46_110,r46_111,r46_112,
		r46_113,r46_114,r46_115,r46_116,r46_117,r46_118,r46_119,r46_120,r46_121,r46_122,r46_123,r46_124,r46_125,r46_126,
	r47_0,r47_1,r47_2,r47_3,r47_4,r47_5,r47_6,r47_7,r47_8,r47_9,r47_10,r47_11,r47_12,r47_13,r47_14,r47_15,r47_16,
		r47_17,r47_18,r47_19,r47_20,r47_21,r47_22,r47_23,r47_24,r47_25,r47_26,r47_27,r47_28,r47_29,r47_30,r47_31,r47_32,
		r47_33,r47_34,r47_35,r47_36,r47_37,r47_38,r47_39,r47_40,r47_41,r47_42,r47_43,r47_44,r47_45,r47_46,r47_47,r47_48,
		r47_49,r47_50,r47_51,r47_52,r47_53,r47_54,r47_55,r47_56,r47_57,r47_58,r47_59,r47_60,r47_61,r47_62,r47_63,r47_64,
		r47_65,r47_66,r47_67,r47_68,r47_69,r47_70,r47_71,r47_72,r47_73,r47_74,r47_75,r47_76,r47_77,r47_78,r47_79,r47_80,
		r47_81,r47_82,r47_83,r47_84,r47_85,r47_86,r47_87,r47_88,r47_89,r47_90,r47_91,r47_92,r47_93,r47_94,r47_95,r47_96,
		r47_97,r47_98,r47_99,r47_100,r47_101,r47_102,r47_103,r47_104,r47_105,r47_106,r47_107,r47_108,r47_109,r47_110,r47_111,r47_112,
		r47_113,r47_114,r47_115,r47_116,r47_117,r47_118,r47_119,r47_120,r47_121,r47_122,r47_123,r47_124,r47_125,r47_126,
	r48_0,r48_1,r48_2,r48_3,r48_4,r48_5,r48_6,r48_7,r48_8,r48_9,r48_10,r48_11,r48_12,r48_13,r48_14,r48_15,r48_16,
		r48_17,r48_18,r48_19,r48_20,r48_21,r48_22,r48_23,r48_24,r48_25,r48_26,r48_27,r48_28,r48_29,r48_30,r48_31,r48_32,
		r48_33,r48_34,r48_35,r48_36,r48_37,r48_38,r48_39,r48_40,r48_41,r48_42,r48_43,r48_44,r48_45,r48_46,r48_47,r48_48,
		r48_49,r48_50,r48_51,r48_52,r48_53,r48_54,r48_55,r48_56,r48_57,r48_58,r48_59,r48_60,r48_61,r48_62,r48_63,r48_64,
		r48_65,r48_66,r48_67,r48_68,r48_69,r48_70,r48_71,r48_72,r48_73,r48_74,r48_75,r48_76,r48_77,r48_78,r48_79,r48_80,
		r48_81,r48_82,r48_83,r48_84,r48_85,r48_86,r48_87,r48_88,r48_89,r48_90,r48_91,r48_92,r48_93,r48_94,r48_95,r48_96,
		r48_97,r48_98,r48_99,r48_100,r48_101,r48_102,r48_103,r48_104,r48_105,r48_106,r48_107,r48_108,r48_109,r48_110,r48_111,r48_112,
		r48_113,r48_114,r48_115,r48_116,r48_117,r48_118,r48_119,r48_120,r48_121,r48_122,r48_123,r48_124,r48_125,r48_126,
	r49_0,r49_1,r49_2,r49_3,r49_4,r49_5,r49_6,r49_7,r49_8,r49_9,r49_10,r49_11,r49_12,r49_13,r49_14,r49_15,r49_16,
		r49_17,r49_18,r49_19,r49_20,r49_21,r49_22,r49_23,r49_24,r49_25,r49_26,r49_27,r49_28,r49_29,r49_30,r49_31,r49_32,
		r49_33,r49_34,r49_35,r49_36,r49_37,r49_38,r49_39,r49_40,r49_41,r49_42,r49_43,r49_44,r49_45,r49_46,r49_47,r49_48,
		r49_49,r49_50,r49_51,r49_52,r49_53,r49_54,r49_55,r49_56,r49_57,r49_58,r49_59,r49_60,r49_61,r49_62,r49_63,r49_64,
		r49_65,r49_66,r49_67,r49_68,r49_69,r49_70,r49_71,r49_72,r49_73,r49_74,r49_75,r49_76,r49_77,r49_78,r49_79,r49_80,
		r49_81,r49_82,r49_83,r49_84,r49_85,r49_86,r49_87,r49_88,r49_89,r49_90,r49_91,r49_92,r49_93,r49_94,r49_95,r49_96,
		r49_97,r49_98,r49_99,r49_100,r49_101,r49_102,r49_103,r49_104,r49_105,r49_106,r49_107,r49_108,r49_109,r49_110,r49_111,r49_112,
		r49_113,r49_114,r49_115,r49_116,r49_117,r49_118,r49_119,r49_120,r49_121,r49_122,r49_123,r49_124,r49_125,r49_126,
	r50_0,r50_1,r50_2,r50_3,r50_4,r50_5,r50_6,r50_7,r50_8,r50_9,r50_10,r50_11,r50_12,r50_13,r50_14,r50_15,r50_16,
		r50_17,r50_18,r50_19,r50_20,r50_21,r50_22,r50_23,r50_24,r50_25,r50_26,r50_27,r50_28,r50_29,r50_30,r50_31,r50_32,
		r50_33,r50_34,r50_35,r50_36,r50_37,r50_38,r50_39,r50_40,r50_41,r50_42,r50_43,r50_44,r50_45,r50_46,r50_47,r50_48,
		r50_49,r50_50,r50_51,r50_52,r50_53,r50_54,r50_55,r50_56,r50_57,r50_58,r50_59,r50_60,r50_61,r50_62,r50_63,r50_64,
		r50_65,r50_66,r50_67,r50_68,r50_69,r50_70,r50_71,r50_72,r50_73,r50_74,r50_75,r50_76,r50_77,r50_78,r50_79,r50_80,
		r50_81,r50_82,r50_83,r50_84,r50_85,r50_86,r50_87,r50_88,r50_89,r50_90,r50_91,r50_92,r50_93,r50_94,r50_95,r50_96,
		r50_97,r50_98,r50_99,r50_100,r50_101,r50_102,r50_103,r50_104,r50_105,r50_106,r50_107,r50_108,r50_109,r50_110,r50_111,r50_112,
		r50_113,r50_114,r50_115,r50_116,r50_117,r50_118,r50_119,r50_120,r50_121,r50_122,r50_123,r50_124,r50_125,r50_126,
	r51_0,r51_1,r51_2,r51_3,r51_4,r51_5,r51_6,r51_7,r51_8,r51_9,r51_10,r51_11,r51_12,r51_13,r51_14,r51_15,r51_16,
		r51_17,r51_18,r51_19,r51_20,r51_21,r51_22,r51_23,r51_24,r51_25,r51_26,r51_27,r51_28,r51_29,r51_30,r51_31,r51_32,
		r51_33,r51_34,r51_35,r51_36,r51_37,r51_38,r51_39,r51_40,r51_41,r51_42,r51_43,r51_44,r51_45,r51_46,r51_47,r51_48,
		r51_49,r51_50,r51_51,r51_52,r51_53,r51_54,r51_55,r51_56,r51_57,r51_58,r51_59,r51_60,r51_61,r51_62,r51_63,r51_64,
		r51_65,r51_66,r51_67,r51_68,r51_69,r51_70,r51_71,r51_72,r51_73,r51_74,r51_75,r51_76,r51_77,r51_78,r51_79,r51_80,
		r51_81,r51_82,r51_83,r51_84,r51_85,r51_86,r51_87,r51_88,r51_89,r51_90,r51_91,r51_92,r51_93,r51_94,r51_95,r51_96,
		r51_97,r51_98,r51_99,r51_100,r51_101,r51_102,r51_103,r51_104,r51_105,r51_106,r51_107,r51_108,r51_109,r51_110,r51_111,r51_112,
		r51_113,r51_114,r51_115,r51_116,r51_117,r51_118,r51_119,r51_120,r51_121,r51_122,r51_123,r51_124,r51_125,r51_126,
	r52_0,r52_1,r52_2,r52_3,r52_4,r52_5,r52_6,r52_7,r52_8,r52_9,r52_10,r52_11,r52_12,r52_13,r52_14,r52_15,r52_16,
		r52_17,r52_18,r52_19,r52_20,r52_21,r52_22,r52_23,r52_24,r52_25,r52_26,r52_27,r52_28,r52_29,r52_30,r52_31,r52_32,
		r52_33,r52_34,r52_35,r52_36,r52_37,r52_38,r52_39,r52_40,r52_41,r52_42,r52_43,r52_44,r52_45,r52_46,r52_47,r52_48,
		r52_49,r52_50,r52_51,r52_52,r52_53,r52_54,r52_55,r52_56,r52_57,r52_58,r52_59,r52_60,r52_61,r52_62,r52_63,r52_64,
		r52_65,r52_66,r52_67,r52_68,r52_69,r52_70,r52_71,r52_72,r52_73,r52_74,r52_75,r52_76,r52_77,r52_78,r52_79,r52_80,
		r52_81,r52_82,r52_83,r52_84,r52_85,r52_86,r52_87,r52_88,r52_89,r52_90,r52_91,r52_92,r52_93,r52_94,r52_95,r52_96,
		r52_97,r52_98,r52_99,r52_100,r52_101,r52_102,r52_103,r52_104,r52_105,r52_106,r52_107,r52_108,r52_109,r52_110,r52_111,r52_112,
		r52_113,r52_114,r52_115,r52_116,r52_117,r52_118,r52_119,r52_120,r52_121,r52_122,r52_123,r52_124,r52_125,r52_126,
	r53_0,r53_1,r53_2,r53_3,r53_4,r53_5,r53_6,r53_7,r53_8,r53_9,r53_10,r53_11,r53_12,r53_13,r53_14,r53_15,r53_16,
		r53_17,r53_18,r53_19,r53_20,r53_21,r53_22,r53_23,r53_24,r53_25,r53_26,r53_27,r53_28,r53_29,r53_30,r53_31,r53_32,
		r53_33,r53_34,r53_35,r53_36,r53_37,r53_38,r53_39,r53_40,r53_41,r53_42,r53_43,r53_44,r53_45,r53_46,r53_47,r53_48,
		r53_49,r53_50,r53_51,r53_52,r53_53,r53_54,r53_55,r53_56,r53_57,r53_58,r53_59,r53_60,r53_61,r53_62,r53_63,r53_64,
		r53_65,r53_66,r53_67,r53_68,r53_69,r53_70,r53_71,r53_72,r53_73,r53_74,r53_75,r53_76,r53_77,r53_78,r53_79,r53_80,
		r53_81,r53_82,r53_83,r53_84,r53_85,r53_86,r53_87,r53_88,r53_89,r53_90,r53_91,r53_92,r53_93,r53_94,r53_95,r53_96,
		r53_97,r53_98,r53_99,r53_100,r53_101,r53_102,r53_103,r53_104,r53_105,r53_106,r53_107,r53_108,r53_109,r53_110,r53_111,r53_112,
		r53_113,r53_114,r53_115,r53_116,r53_117,r53_118,r53_119,r53_120,r53_121,r53_122,r53_123,r53_124,r53_125,r53_126,
	r54_0,r54_1,r54_2,r54_3,r54_4,r54_5,r54_6,r54_7,r54_8,r54_9,r54_10,r54_11,r54_12,r54_13,r54_14,r54_15,r54_16,
		r54_17,r54_18,r54_19,r54_20,r54_21,r54_22,r54_23,r54_24,r54_25,r54_26,r54_27,r54_28,r54_29,r54_30,r54_31,r54_32,
		r54_33,r54_34,r54_35,r54_36,r54_37,r54_38,r54_39,r54_40,r54_41,r54_42,r54_43,r54_44,r54_45,r54_46,r54_47,r54_48,
		r54_49,r54_50,r54_51,r54_52,r54_53,r54_54,r54_55,r54_56,r54_57,r54_58,r54_59,r54_60,r54_61,r54_62,r54_63,r54_64,
		r54_65,r54_66,r54_67,r54_68,r54_69,r54_70,r54_71,r54_72,r54_73,r54_74,r54_75,r54_76,r54_77,r54_78,r54_79,r54_80,
		r54_81,r54_82,r54_83,r54_84,r54_85,r54_86,r54_87,r54_88,r54_89,r54_90,r54_91,r54_92,r54_93,r54_94,r54_95,r54_96,
		r54_97,r54_98,r54_99,r54_100,r54_101,r54_102,r54_103,r54_104,r54_105,r54_106,r54_107,r54_108,r54_109,r54_110,r54_111,r54_112,
		r54_113,r54_114,r54_115,r54_116,r54_117,r54_118,r54_119,r54_120,r54_121,r54_122,r54_123,r54_124,r54_125,r54_126,
	r55_0,r55_1,r55_2,r55_3,r55_4,r55_5,r55_6,r55_7,r55_8,r55_9,r55_10,r55_11,r55_12,r55_13,r55_14,r55_15,r55_16,
		r55_17,r55_18,r55_19,r55_20,r55_21,r55_22,r55_23,r55_24,r55_25,r55_26,r55_27,r55_28,r55_29,r55_30,r55_31,r55_32,
		r55_33,r55_34,r55_35,r55_36,r55_37,r55_38,r55_39,r55_40,r55_41,r55_42,r55_43,r55_44,r55_45,r55_46,r55_47,r55_48,
		r55_49,r55_50,r55_51,r55_52,r55_53,r55_54,r55_55,r55_56,r55_57,r55_58,r55_59,r55_60,r55_61,r55_62,r55_63,r55_64,
		r55_65,r55_66,r55_67,r55_68,r55_69,r55_70,r55_71,r55_72,r55_73,r55_74,r55_75,r55_76,r55_77,r55_78,r55_79,r55_80,
		r55_81,r55_82,r55_83,r55_84,r55_85,r55_86,r55_87,r55_88,r55_89,r55_90,r55_91,r55_92,r55_93,r55_94,r55_95,r55_96,
		r55_97,r55_98,r55_99,r55_100,r55_101,r55_102,r55_103,r55_104,r55_105,r55_106,r55_107,r55_108,r55_109,r55_110,r55_111,r55_112,
		r55_113,r55_114,r55_115,r55_116,r55_117,r55_118,r55_119,r55_120,r55_121,r55_122,r55_123,r55_124,r55_125,r55_126,
	r56_0,r56_1,r56_2,r56_3,r56_4,r56_5,r56_6,r56_7,r56_8,r56_9,r56_10,r56_11,r56_12,r56_13,r56_14,r56_15,r56_16,
		r56_17,r56_18,r56_19,r56_20,r56_21,r56_22,r56_23,r56_24,r56_25,r56_26,r56_27,r56_28,r56_29,r56_30,r56_31,r56_32,
		r56_33,r56_34,r56_35,r56_36,r56_37,r56_38,r56_39,r56_40,r56_41,r56_42,r56_43,r56_44,r56_45,r56_46,r56_47,r56_48,
		r56_49,r56_50,r56_51,r56_52,r56_53,r56_54,r56_55,r56_56,r56_57,r56_58,r56_59,r56_60,r56_61,r56_62,r56_63,r56_64,
		r56_65,r56_66,r56_67,r56_68,r56_69,r56_70,r56_71,r56_72,r56_73,r56_74,r56_75,r56_76,r56_77,r56_78,r56_79,r56_80,
		r56_81,r56_82,r56_83,r56_84,r56_85,r56_86,r56_87,r56_88,r56_89,r56_90,r56_91,r56_92,r56_93,r56_94,r56_95,r56_96,
		r56_97,r56_98,r56_99,r56_100,r56_101,r56_102,r56_103,r56_104,r56_105,r56_106,r56_107,r56_108,r56_109,r56_110,r56_111,r56_112,
		r56_113,r56_114,r56_115,r56_116,r56_117,r56_118,r56_119,r56_120,r56_121,r56_122,r56_123,r56_124,r56_125,r56_126,
	r57_0,r57_1,r57_2,r57_3,r57_4,r57_5,r57_6,r57_7,r57_8,r57_9,r57_10,r57_11,r57_12,r57_13,r57_14,r57_15,r57_16,
		r57_17,r57_18,r57_19,r57_20,r57_21,r57_22,r57_23,r57_24,r57_25,r57_26,r57_27,r57_28,r57_29,r57_30,r57_31,r57_32,
		r57_33,r57_34,r57_35,r57_36,r57_37,r57_38,r57_39,r57_40,r57_41,r57_42,r57_43,r57_44,r57_45,r57_46,r57_47,r57_48,
		r57_49,r57_50,r57_51,r57_52,r57_53,r57_54,r57_55,r57_56,r57_57,r57_58,r57_59,r57_60,r57_61,r57_62,r57_63,r57_64,
		r57_65,r57_66,r57_67,r57_68,r57_69,r57_70,r57_71,r57_72,r57_73,r57_74,r57_75,r57_76,r57_77,r57_78,r57_79,r57_80,
		r57_81,r57_82,r57_83,r57_84,r57_85,r57_86,r57_87,r57_88,r57_89,r57_90,r57_91,r57_92,r57_93,r57_94,r57_95,r57_96,
		r57_97,r57_98,r57_99,r57_100,r57_101,r57_102,r57_103,r57_104,r57_105,r57_106,r57_107,r57_108,r57_109,r57_110,r57_111,r57_112,
		r57_113,r57_114,r57_115,r57_116,r57_117,r57_118,r57_119,r57_120,r57_121,r57_122,r57_123,r57_124,r57_125,r57_126,
	r58_0,r58_1,r58_2,r58_3,r58_4,r58_5,r58_6,r58_7,r58_8,r58_9,r58_10,r58_11,r58_12,r58_13,r58_14,r58_15,r58_16,
		r58_17,r58_18,r58_19,r58_20,r58_21,r58_22,r58_23,r58_24,r58_25,r58_26,r58_27,r58_28,r58_29,r58_30,r58_31,r58_32,
		r58_33,r58_34,r58_35,r58_36,r58_37,r58_38,r58_39,r58_40,r58_41,r58_42,r58_43,r58_44,r58_45,r58_46,r58_47,r58_48,
		r58_49,r58_50,r58_51,r58_52,r58_53,r58_54,r58_55,r58_56,r58_57,r58_58,r58_59,r58_60,r58_61,r58_62,r58_63,r58_64,
		r58_65,r58_66,r58_67,r58_68,r58_69,r58_70,r58_71,r58_72,r58_73,r58_74,r58_75,r58_76,r58_77,r58_78,r58_79,r58_80,
		r58_81,r58_82,r58_83,r58_84,r58_85,r58_86,r58_87,r58_88,r58_89,r58_90,r58_91,r58_92,r58_93,r58_94,r58_95,r58_96,
		r58_97,r58_98,r58_99,r58_100,r58_101,r58_102,r58_103,r58_104,r58_105,r58_106,r58_107,r58_108,r58_109,r58_110,r58_111,r58_112,
		r58_113,r58_114,r58_115,r58_116,r58_117,r58_118,r58_119,r58_120,r58_121,r58_122,r58_123,r58_124,r58_125,r58_126,
	r59_0,r59_1,r59_2,r59_3,r59_4,r59_5,r59_6,r59_7,r59_8,r59_9,r59_10,r59_11,r59_12,r59_13,r59_14,r59_15,r59_16,
		r59_17,r59_18,r59_19,r59_20,r59_21,r59_22,r59_23,r59_24,r59_25,r59_26,r59_27,r59_28,r59_29,r59_30,r59_31,r59_32,
		r59_33,r59_34,r59_35,r59_36,r59_37,r59_38,r59_39,r59_40,r59_41,r59_42,r59_43,r59_44,r59_45,r59_46,r59_47,r59_48,
		r59_49,r59_50,r59_51,r59_52,r59_53,r59_54,r59_55,r59_56,r59_57,r59_58,r59_59,r59_60,r59_61,r59_62,r59_63,r59_64,
		r59_65,r59_66,r59_67,r59_68,r59_69,r59_70,r59_71,r59_72,r59_73,r59_74,r59_75,r59_76,r59_77,r59_78,r59_79,r59_80,
		r59_81,r59_82,r59_83,r59_84,r59_85,r59_86,r59_87,r59_88,r59_89,r59_90,r59_91,r59_92,r59_93,r59_94,r59_95,r59_96,
		r59_97,r59_98,r59_99,r59_100,r59_101,r59_102,r59_103,r59_104,r59_105,r59_106,r59_107,r59_108,r59_109,r59_110,r59_111,r59_112,
		r59_113,r59_114,r59_115,r59_116,r59_117,r59_118,r59_119,r59_120,r59_121,r59_122,r59_123,r59_124,r59_125,r59_126,
	r60_0,r60_1,r60_2,r60_3,r60_4,r60_5,r60_6,r60_7,r60_8,r60_9,r60_10,r60_11,r60_12,r60_13,r60_14,r60_15,r60_16,
		r60_17,r60_18,r60_19,r60_20,r60_21,r60_22,r60_23,r60_24,r60_25,r60_26,r60_27,r60_28,r60_29,r60_30,r60_31,r60_32,
		r60_33,r60_34,r60_35,r60_36,r60_37,r60_38,r60_39,r60_40,r60_41,r60_42,r60_43,r60_44,r60_45,r60_46,r60_47,r60_48,
		r60_49,r60_50,r60_51,r60_52,r60_53,r60_54,r60_55,r60_56,r60_57,r60_58,r60_59,r60_60,r60_61,r60_62,r60_63,r60_64,
		r60_65,r60_66,r60_67,r60_68,r60_69,r60_70,r60_71,r60_72,r60_73,r60_74,r60_75,r60_76,r60_77,r60_78,r60_79,r60_80,
		r60_81,r60_82,r60_83,r60_84,r60_85,r60_86,r60_87,r60_88,r60_89,r60_90,r60_91,r60_92,r60_93,r60_94,r60_95,r60_96,
		r60_97,r60_98,r60_99,r60_100,r60_101,r60_102,r60_103,r60_104,r60_105,r60_106,r60_107,r60_108,r60_109,r60_110,r60_111,r60_112,
		r60_113,r60_114,r60_115,r60_116,r60_117,r60_118,r60_119,r60_120,r60_121,r60_122,r60_123,r60_124,r60_125,r60_126,
	r61_0,r61_1,r61_2,r61_3,r61_4,r61_5,r61_6,r61_7,r61_8,r61_9,r61_10,r61_11,r61_12,r61_13,r61_14,r61_15,r61_16,
		r61_17,r61_18,r61_19,r61_20,r61_21,r61_22,r61_23,r61_24,r61_25,r61_26,r61_27,r61_28,r61_29,r61_30,r61_31,r61_32,
		r61_33,r61_34,r61_35,r61_36,r61_37,r61_38,r61_39,r61_40,r61_41,r61_42,r61_43,r61_44,r61_45,r61_46,r61_47,r61_48,
		r61_49,r61_50,r61_51,r61_52,r61_53,r61_54,r61_55,r61_56,r61_57,r61_58,r61_59,r61_60,r61_61,r61_62,r61_63,r61_64,
		r61_65,r61_66,r61_67,r61_68,r61_69,r61_70,r61_71,r61_72,r61_73,r61_74,r61_75,r61_76,r61_77,r61_78,r61_79,r61_80,
		r61_81,r61_82,r61_83,r61_84,r61_85,r61_86,r61_87,r61_88,r61_89,r61_90,r61_91,r61_92,r61_93,r61_94,r61_95,r61_96,
		r61_97,r61_98,r61_99,r61_100,r61_101,r61_102,r61_103,r61_104,r61_105,r61_106,r61_107,r61_108,r61_109,r61_110,r61_111,r61_112,
		r61_113,r61_114,r61_115,r61_116,r61_117,r61_118,r61_119,r61_120,r61_121,r61_122,r61_123,r61_124,r61_125,r61_126,
	r62_0,r62_1,r62_2,r62_3,r62_4,r62_5,r62_6,r62_7,r62_8,r62_9,r62_10,r62_11,r62_12,r62_13,r62_14,r62_15,r62_16,
		r62_17,r62_18,r62_19,r62_20,r62_21,r62_22,r62_23,r62_24,r62_25,r62_26,r62_27,r62_28,r62_29,r62_30,r62_31,r62_32,
		r62_33,r62_34,r62_35,r62_36,r62_37,r62_38,r62_39,r62_40,r62_41,r62_42,r62_43,r62_44,r62_45,r62_46,r62_47,r62_48,
		r62_49,r62_50,r62_51,r62_52,r62_53,r62_54,r62_55,r62_56,r62_57,r62_58,r62_59,r62_60,r62_61,r62_62,r62_63,r62_64,
		r62_65,r62_66,r62_67,r62_68,r62_69,r62_70,r62_71,r62_72,r62_73,r62_74,r62_75,r62_76,r62_77,r62_78,r62_79,r62_80,
		r62_81,r62_82,r62_83,r62_84,r62_85,r62_86,r62_87,r62_88,r62_89,r62_90,r62_91,r62_92,r62_93,r62_94,r62_95,r62_96,
		r62_97,r62_98,r62_99,r62_100,r62_101,r62_102,r62_103,r62_104,r62_105,r62_106,r62_107,r62_108,r62_109,r62_110,r62_111,r62_112,
		r62_113,r62_114,r62_115,r62_116,r62_117,r62_118,r62_119,r62_120,r62_121,r62_122,r62_123,r62_124,r62_125,r62_126,
	r63_0,r63_1,r63_2,r63_3,r63_4,r63_5,r63_6,r63_7,r63_8,r63_9,r63_10,r63_11,r63_12,r63_13,r63_14,r63_15,r63_16,
		r63_17,r63_18,r63_19,r63_20,r63_21,r63_22,r63_23,r63_24,r63_25,r63_26,r63_27,r63_28,r63_29,r63_30,r63_31,r63_32,
		r63_33,r63_34,r63_35,r63_36,r63_37,r63_38,r63_39,r63_40,r63_41,r63_42,r63_43,r63_44,r63_45,r63_46,r63_47,r63_48,
		r63_49,r63_50,r63_51,r63_52,r63_53,r63_54,r63_55,r63_56,r63_57,r63_58,r63_59,r63_60,r63_61,r63_62,r63_63,r63_64,
		r63_65,r63_66,r63_67,r63_68,r63_69,r63_70,r63_71,r63_72,r63_73,r63_74,r63_75,r63_76,r63_77,r63_78,r63_79,r63_80,
		r63_81,r63_82,r63_83,r63_84,r63_85,r63_86,r63_87,r63_88,r63_89,r63_90,r63_91,r63_92,r63_93,r63_94,r63_95,r63_96,
		r63_97,r63_98,r63_99,r63_100,r63_101,r63_102,r63_103,r63_104,r63_105,r63_106,r63_107,r63_108,r63_109,r63_110,r63_111,r63_112,
		r63_113,r63_114,r63_115,r63_116,r63_117,r63_118,r63_119,r63_120,r63_121,r63_122,r63_123,r63_124,r63_125,r63_126,
	r64_0,r64_1,r64_2,r64_3,r64_4,r64_5,r64_6,r64_7,r64_8,r64_9,r64_10,r64_11,r64_12,r64_13,r64_14,r64_15,r64_16,
		r64_17,r64_18,r64_19,r64_20,r64_21,r64_22,r64_23,r64_24,r64_25,r64_26,r64_27,r64_28,r64_29,r64_30,r64_31,r64_32,
		r64_33,r64_34,r64_35,r64_36,r64_37,r64_38,r64_39,r64_40,r64_41,r64_42,r64_43,r64_44,r64_45,r64_46,r64_47,r64_48,
		r64_49,r64_50,r64_51,r64_52,r64_53,r64_54,r64_55,r64_56,r64_57,r64_58,r64_59,r64_60,r64_61,r64_62,r64_63,r64_64,
		r64_65,r64_66,r64_67,r64_68,r64_69,r64_70,r64_71,r64_72,r64_73,r64_74,r64_75,r64_76,r64_77,r64_78,r64_79,r64_80,
		r64_81,r64_82,r64_83,r64_84,r64_85,r64_86,r64_87,r64_88,r64_89,r64_90,r64_91,r64_92,r64_93,r64_94,r64_95,r64_96,
		r64_97,r64_98,r64_99,r64_100,r64_101,r64_102,r64_103,r64_104,r64_105,r64_106,r64_107,r64_108,r64_109,r64_110,r64_111,r64_112,
		r64_113,r64_114,r64_115,r64_116,r64_117,r64_118,r64_119,r64_120,r64_121,r64_122,r64_123,r64_124,r64_125,r64_126,
	r65_0,r65_1,r65_2,r65_3,r65_4,r65_5,r65_6,r65_7,r65_8,r65_9,r65_10,r65_11,r65_12,r65_13,r65_14,r65_15,r65_16,
		r65_17,r65_18,r65_19,r65_20,r65_21,r65_22,r65_23,r65_24,r65_25,r65_26,r65_27,r65_28,r65_29,r65_30,r65_31,r65_32,
		r65_33,r65_34,r65_35,r65_36,r65_37,r65_38,r65_39,r65_40,r65_41,r65_42,r65_43,r65_44,r65_45,r65_46,r65_47,r65_48,
		r65_49,r65_50,r65_51,r65_52,r65_53,r65_54,r65_55,r65_56,r65_57,r65_58,r65_59,r65_60,r65_61,r65_62,r65_63,r65_64,
		r65_65,r65_66,r65_67,r65_68,r65_69,r65_70,r65_71,r65_72,r65_73,r65_74,r65_75,r65_76,r65_77,r65_78,r65_79,r65_80,
		r65_81,r65_82,r65_83,r65_84,r65_85,r65_86,r65_87,r65_88,r65_89,r65_90,r65_91,r65_92,r65_93,r65_94,r65_95,r65_96,
		r65_97,r65_98,r65_99,r65_100,r65_101,r65_102,r65_103,r65_104,r65_105,r65_106,r65_107,r65_108,r65_109,r65_110,r65_111,r65_112,
		r65_113,r65_114,r65_115,r65_116,r65_117,r65_118,r65_119,r65_120,r65_121,r65_122,r65_123,r65_124,r65_125,r65_126,
	r66_0,r66_1,r66_2,r66_3,r66_4,r66_5,r66_6,r66_7,r66_8,r66_9,r66_10,r66_11,r66_12,r66_13,r66_14,r66_15,r66_16,
		r66_17,r66_18,r66_19,r66_20,r66_21,r66_22,r66_23,r66_24,r66_25,r66_26,r66_27,r66_28,r66_29,r66_30,r66_31,r66_32,
		r66_33,r66_34,r66_35,r66_36,r66_37,r66_38,r66_39,r66_40,r66_41,r66_42,r66_43,r66_44,r66_45,r66_46,r66_47,r66_48,
		r66_49,r66_50,r66_51,r66_52,r66_53,r66_54,r66_55,r66_56,r66_57,r66_58,r66_59,r66_60,r66_61,r66_62,r66_63,r66_64,
		r66_65,r66_66,r66_67,r66_68,r66_69,r66_70,r66_71,r66_72,r66_73,r66_74,r66_75,r66_76,r66_77,r66_78,r66_79,r66_80,
		r66_81,r66_82,r66_83,r66_84,r66_85,r66_86,r66_87,r66_88,r66_89,r66_90,r66_91,r66_92,r66_93,r66_94,r66_95,r66_96,
		r66_97,r66_98,r66_99,r66_100,r66_101,r66_102,r66_103,r66_104,r66_105,r66_106,r66_107,r66_108,r66_109,r66_110,r66_111,r66_112,
		r66_113,r66_114,r66_115,r66_116,r66_117,r66_118,r66_119,r66_120,r66_121,r66_122,r66_123,r66_124,r66_125,r66_126,
	r67_0,r67_1,r67_2,r67_3,r67_4,r67_5,r67_6,r67_7,r67_8,r67_9,r67_10,r67_11,r67_12,r67_13,r67_14,r67_15,r67_16,
		r67_17,r67_18,r67_19,r67_20,r67_21,r67_22,r67_23,r67_24,r67_25,r67_26,r67_27,r67_28,r67_29,r67_30,r67_31,r67_32,
		r67_33,r67_34,r67_35,r67_36,r67_37,r67_38,r67_39,r67_40,r67_41,r67_42,r67_43,r67_44,r67_45,r67_46,r67_47,r67_48,
		r67_49,r67_50,r67_51,r67_52,r67_53,r67_54,r67_55,r67_56,r67_57,r67_58,r67_59,r67_60,r67_61,r67_62,r67_63,r67_64,
		r67_65,r67_66,r67_67,r67_68,r67_69,r67_70,r67_71,r67_72,r67_73,r67_74,r67_75,r67_76,r67_77,r67_78,r67_79,r67_80,
		r67_81,r67_82,r67_83,r67_84,r67_85,r67_86,r67_87,r67_88,r67_89,r67_90,r67_91,r67_92,r67_93,r67_94,r67_95,r67_96,
		r67_97,r67_98,r67_99,r67_100,r67_101,r67_102,r67_103,r67_104,r67_105,r67_106,r67_107,r67_108,r67_109,r67_110,r67_111,r67_112,
		r67_113,r67_114,r67_115,r67_116,r67_117,r67_118,r67_119,r67_120,r67_121,r67_122,r67_123,r67_124,r67_125,r67_126,
	r68_0,r68_1,r68_2,r68_3,r68_4,r68_5,r68_6,r68_7,r68_8,r68_9,r68_10,r68_11,r68_12,r68_13,r68_14,r68_15,r68_16,
		r68_17,r68_18,r68_19,r68_20,r68_21,r68_22,r68_23,r68_24,r68_25,r68_26,r68_27,r68_28,r68_29,r68_30,r68_31,r68_32,
		r68_33,r68_34,r68_35,r68_36,r68_37,r68_38,r68_39,r68_40,r68_41,r68_42,r68_43,r68_44,r68_45,r68_46,r68_47,r68_48,
		r68_49,r68_50,r68_51,r68_52,r68_53,r68_54,r68_55,r68_56,r68_57,r68_58,r68_59,r68_60,r68_61,r68_62,r68_63,r68_64,
		r68_65,r68_66,r68_67,r68_68,r68_69,r68_70,r68_71,r68_72,r68_73,r68_74,r68_75,r68_76,r68_77,r68_78,r68_79,r68_80,
		r68_81,r68_82,r68_83,r68_84,r68_85,r68_86,r68_87,r68_88,r68_89,r68_90,r68_91,r68_92,r68_93,r68_94,r68_95,r68_96,
		r68_97,r68_98,r68_99,r68_100,r68_101,r68_102,r68_103,r68_104,r68_105,r68_106,r68_107,r68_108,r68_109,r68_110,r68_111,r68_112,
		r68_113,r68_114,r68_115,r68_116,r68_117,r68_118,r68_119,r68_120,r68_121,r68_122,r68_123,r68_124,r68_125,r68_126,
	r69_0,r69_1,r69_2,r69_3,r69_4,r69_5,r69_6,r69_7,r69_8,r69_9,r69_10,r69_11,r69_12,r69_13,r69_14,r69_15,r69_16,
		r69_17,r69_18,r69_19,r69_20,r69_21,r69_22,r69_23,r69_24,r69_25,r69_26,r69_27,r69_28,r69_29,r69_30,r69_31,r69_32,
		r69_33,r69_34,r69_35,r69_36,r69_37,r69_38,r69_39,r69_40,r69_41,r69_42,r69_43,r69_44,r69_45,r69_46,r69_47,r69_48,
		r69_49,r69_50,r69_51,r69_52,r69_53,r69_54,r69_55,r69_56,r69_57,r69_58,r69_59,r69_60,r69_61,r69_62,r69_63,r69_64,
		r69_65,r69_66,r69_67,r69_68,r69_69,r69_70,r69_71,r69_72,r69_73,r69_74,r69_75,r69_76,r69_77,r69_78,r69_79,r69_80,
		r69_81,r69_82,r69_83,r69_84,r69_85,r69_86,r69_87,r69_88,r69_89,r69_90,r69_91,r69_92,r69_93,r69_94,r69_95,r69_96,
		r69_97,r69_98,r69_99,r69_100,r69_101,r69_102,r69_103,r69_104,r69_105,r69_106,r69_107,r69_108,r69_109,r69_110,r69_111,r69_112,
		r69_113,r69_114,r69_115,r69_116,r69_117,r69_118,r69_119,r69_120,r69_121,r69_122,r69_123,r69_124,r69_125,r69_126,
	r70_0,r70_1,r70_2,r70_3,r70_4,r70_5,r70_6,r70_7,r70_8,r70_9,r70_10,r70_11,r70_12,r70_13,r70_14,r70_15,r70_16,
		r70_17,r70_18,r70_19,r70_20,r70_21,r70_22,r70_23,r70_24,r70_25,r70_26,r70_27,r70_28,r70_29,r70_30,r70_31,r70_32,
		r70_33,r70_34,r70_35,r70_36,r70_37,r70_38,r70_39,r70_40,r70_41,r70_42,r70_43,r70_44,r70_45,r70_46,r70_47,r70_48,
		r70_49,r70_50,r70_51,r70_52,r70_53,r70_54,r70_55,r70_56,r70_57,r70_58,r70_59,r70_60,r70_61,r70_62,r70_63,r70_64,
		r70_65,r70_66,r70_67,r70_68,r70_69,r70_70,r70_71,r70_72,r70_73,r70_74,r70_75,r70_76,r70_77,r70_78,r70_79,r70_80,
		r70_81,r70_82,r70_83,r70_84,r70_85,r70_86,r70_87,r70_88,r70_89,r70_90,r70_91,r70_92,r70_93,r70_94,r70_95,r70_96,
		r70_97,r70_98,r70_99,r70_100,r70_101,r70_102,r70_103,r70_104,r70_105,r70_106,r70_107,r70_108,r70_109,r70_110,r70_111,r70_112,
		r70_113,r70_114,r70_115,r70_116,r70_117,r70_118,r70_119,r70_120,r70_121,r70_122,r70_123,r70_124,r70_125,r70_126,
	r71_0,r71_1,r71_2,r71_3,r71_4,r71_5,r71_6,r71_7,r71_8,r71_9,r71_10,r71_11,r71_12,r71_13,r71_14,r71_15,r71_16,
		r71_17,r71_18,r71_19,r71_20,r71_21,r71_22,r71_23,r71_24,r71_25,r71_26,r71_27,r71_28,r71_29,r71_30,r71_31,r71_32,
		r71_33,r71_34,r71_35,r71_36,r71_37,r71_38,r71_39,r71_40,r71_41,r71_42,r71_43,r71_44,r71_45,r71_46,r71_47,r71_48,
		r71_49,r71_50,r71_51,r71_52,r71_53,r71_54,r71_55,r71_56,r71_57,r71_58,r71_59,r71_60,r71_61,r71_62,r71_63,r71_64,
		r71_65,r71_66,r71_67,r71_68,r71_69,r71_70,r71_71,r71_72,r71_73,r71_74,r71_75,r71_76,r71_77,r71_78,r71_79,r71_80,
		r71_81,r71_82,r71_83,r71_84,r71_85,r71_86,r71_87,r71_88,r71_89,r71_90,r71_91,r71_92,r71_93,r71_94,r71_95,r71_96,
		r71_97,r71_98,r71_99,r71_100,r71_101,r71_102,r71_103,r71_104,r71_105,r71_106,r71_107,r71_108,r71_109,r71_110,r71_111,r71_112,
		r71_113,r71_114,r71_115,r71_116,r71_117,r71_118,r71_119,r71_120,r71_121,r71_122,r71_123,r71_124,r71_125,r71_126,
	r72_0,r72_1,r72_2,r72_3,r72_4,r72_5,r72_6,r72_7,r72_8,r72_9,r72_10,r72_11,r72_12,r72_13,r72_14,r72_15,r72_16,
		r72_17,r72_18,r72_19,r72_20,r72_21,r72_22,r72_23,r72_24,r72_25,r72_26,r72_27,r72_28,r72_29,r72_30,r72_31,r72_32,
		r72_33,r72_34,r72_35,r72_36,r72_37,r72_38,r72_39,r72_40,r72_41,r72_42,r72_43,r72_44,r72_45,r72_46,r72_47,r72_48,
		r72_49,r72_50,r72_51,r72_52,r72_53,r72_54,r72_55,r72_56,r72_57,r72_58,r72_59,r72_60,r72_61,r72_62,r72_63,r72_64,
		r72_65,r72_66,r72_67,r72_68,r72_69,r72_70,r72_71,r72_72,r72_73,r72_74,r72_75,r72_76,r72_77,r72_78,r72_79,r72_80,
		r72_81,r72_82,r72_83,r72_84,r72_85,r72_86,r72_87,r72_88,r72_89,r72_90,r72_91,r72_92,r72_93,r72_94,r72_95,r72_96,
		r72_97,r72_98,r72_99,r72_100,r72_101,r72_102,r72_103,r72_104,r72_105,r72_106,r72_107,r72_108,r72_109,r72_110,r72_111,r72_112,
		r72_113,r72_114,r72_115,r72_116,r72_117,r72_118,r72_119,r72_120,r72_121,r72_122,r72_123,r72_124,r72_125,r72_126,
	r73_0,r73_1,r73_2,r73_3,r73_4,r73_5,r73_6,r73_7,r73_8,r73_9,r73_10,r73_11,r73_12,r73_13,r73_14,r73_15,r73_16,
		r73_17,r73_18,r73_19,r73_20,r73_21,r73_22,r73_23,r73_24,r73_25,r73_26,r73_27,r73_28,r73_29,r73_30,r73_31,r73_32,
		r73_33,r73_34,r73_35,r73_36,r73_37,r73_38,r73_39,r73_40,r73_41,r73_42,r73_43,r73_44,r73_45,r73_46,r73_47,r73_48,
		r73_49,r73_50,r73_51,r73_52,r73_53,r73_54,r73_55,r73_56,r73_57,r73_58,r73_59,r73_60,r73_61,r73_62,r73_63,r73_64,
		r73_65,r73_66,r73_67,r73_68,r73_69,r73_70,r73_71,r73_72,r73_73,r73_74,r73_75,r73_76,r73_77,r73_78,r73_79,r73_80,
		r73_81,r73_82,r73_83,r73_84,r73_85,r73_86,r73_87,r73_88,r73_89,r73_90,r73_91,r73_92,r73_93,r73_94,r73_95,r73_96,
		r73_97,r73_98,r73_99,r73_100,r73_101,r73_102,r73_103,r73_104,r73_105,r73_106,r73_107,r73_108,r73_109,r73_110,r73_111,r73_112,
		r73_113,r73_114,r73_115,r73_116,r73_117,r73_118,r73_119,r73_120,r73_121,r73_122,r73_123,r73_124,r73_125,r73_126,
	r74_0,r74_1,r74_2,r74_3,r74_4,r74_5,r74_6,r74_7,r74_8,r74_9,r74_10,r74_11,r74_12,r74_13,r74_14,r74_15,r74_16,
		r74_17,r74_18,r74_19,r74_20,r74_21,r74_22,r74_23,r74_24,r74_25,r74_26,r74_27,r74_28,r74_29,r74_30,r74_31,r74_32,
		r74_33,r74_34,r74_35,r74_36,r74_37,r74_38,r74_39,r74_40,r74_41,r74_42,r74_43,r74_44,r74_45,r74_46,r74_47,r74_48,
		r74_49,r74_50,r74_51,r74_52,r74_53,r74_54,r74_55,r74_56,r74_57,r74_58,r74_59,r74_60,r74_61,r74_62,r74_63,r74_64,
		r74_65,r74_66,r74_67,r74_68,r74_69,r74_70,r74_71,r74_72,r74_73,r74_74,r74_75,r74_76,r74_77,r74_78,r74_79,r74_80,
		r74_81,r74_82,r74_83,r74_84,r74_85,r74_86,r74_87,r74_88,r74_89,r74_90,r74_91,r74_92,r74_93,r74_94,r74_95,r74_96,
		r74_97,r74_98,r74_99,r74_100,r74_101,r74_102,r74_103,r74_104,r74_105,r74_106,r74_107,r74_108,r74_109,r74_110,r74_111,r74_112,
		r74_113,r74_114,r74_115,r74_116,r74_117,r74_118,r74_119,r74_120,r74_121,r74_122,r74_123,r74_124,r74_125,r74_126,
	r75_0,r75_1,r75_2,r75_3,r75_4,r75_5,r75_6,r75_7,r75_8,r75_9,r75_10,r75_11,r75_12,r75_13,r75_14,r75_15,r75_16,
		r75_17,r75_18,r75_19,r75_20,r75_21,r75_22,r75_23,r75_24,r75_25,r75_26,r75_27,r75_28,r75_29,r75_30,r75_31,r75_32,
		r75_33,r75_34,r75_35,r75_36,r75_37,r75_38,r75_39,r75_40,r75_41,r75_42,r75_43,r75_44,r75_45,r75_46,r75_47,r75_48,
		r75_49,r75_50,r75_51,r75_52,r75_53,r75_54,r75_55,r75_56,r75_57,r75_58,r75_59,r75_60,r75_61,r75_62,r75_63,r75_64,
		r75_65,r75_66,r75_67,r75_68,r75_69,r75_70,r75_71,r75_72,r75_73,r75_74,r75_75,r75_76,r75_77,r75_78,r75_79,r75_80,
		r75_81,r75_82,r75_83,r75_84,r75_85,r75_86,r75_87,r75_88,r75_89,r75_90,r75_91,r75_92,r75_93,r75_94,r75_95,r75_96,
		r75_97,r75_98,r75_99,r75_100,r75_101,r75_102,r75_103,r75_104,r75_105,r75_106,r75_107,r75_108,r75_109,r75_110,r75_111,r75_112,
		r75_113,r75_114,r75_115,r75_116,r75_117,r75_118,r75_119,r75_120,r75_121,r75_122,r75_123,r75_124,r75_125,r75_126,
	r76_0,r76_1,r76_2,r76_3,r76_4,r76_5,r76_6,r76_7,r76_8,r76_9,r76_10,r76_11,r76_12,r76_13,r76_14,r76_15,r76_16,
		r76_17,r76_18,r76_19,r76_20,r76_21,r76_22,r76_23,r76_24,r76_25,r76_26,r76_27,r76_28,r76_29,r76_30,r76_31,r76_32,
		r76_33,r76_34,r76_35,r76_36,r76_37,r76_38,r76_39,r76_40,r76_41,r76_42,r76_43,r76_44,r76_45,r76_46,r76_47,r76_48,
		r76_49,r76_50,r76_51,r76_52,r76_53,r76_54,r76_55,r76_56,r76_57,r76_58,r76_59,r76_60,r76_61,r76_62,r76_63,r76_64,
		r76_65,r76_66,r76_67,r76_68,r76_69,r76_70,r76_71,r76_72,r76_73,r76_74,r76_75,r76_76,r76_77,r76_78,r76_79,r76_80,
		r76_81,r76_82,r76_83,r76_84,r76_85,r76_86,r76_87,r76_88,r76_89,r76_90,r76_91,r76_92,r76_93,r76_94,r76_95,r76_96,
		r76_97,r76_98,r76_99,r76_100,r76_101,r76_102,r76_103,r76_104,r76_105,r76_106,r76_107,r76_108,r76_109,r76_110,r76_111,r76_112,
		r76_113,r76_114,r76_115,r76_116,r76_117,r76_118,r76_119,r76_120,r76_121,r76_122,r76_123,r76_124,r76_125,r76_126,
	r77_0,r77_1,r77_2,r77_3,r77_4,r77_5,r77_6,r77_7,r77_8,r77_9,r77_10,r77_11,r77_12,r77_13,r77_14,r77_15,r77_16,
		r77_17,r77_18,r77_19,r77_20,r77_21,r77_22,r77_23,r77_24,r77_25,r77_26,r77_27,r77_28,r77_29,r77_30,r77_31,r77_32,
		r77_33,r77_34,r77_35,r77_36,r77_37,r77_38,r77_39,r77_40,r77_41,r77_42,r77_43,r77_44,r77_45,r77_46,r77_47,r77_48,
		r77_49,r77_50,r77_51,r77_52,r77_53,r77_54,r77_55,r77_56,r77_57,r77_58,r77_59,r77_60,r77_61,r77_62,r77_63,r77_64,
		r77_65,r77_66,r77_67,r77_68,r77_69,r77_70,r77_71,r77_72,r77_73,r77_74,r77_75,r77_76,r77_77,r77_78,r77_79,r77_80,
		r77_81,r77_82,r77_83,r77_84,r77_85,r77_86,r77_87,r77_88,r77_89,r77_90,r77_91,r77_92,r77_93,r77_94,r77_95,r77_96,
		r77_97,r77_98,r77_99,r77_100,r77_101,r77_102,r77_103,r77_104,r77_105,r77_106,r77_107,r77_108,r77_109,r77_110,r77_111,r77_112,
		r77_113,r77_114,r77_115,r77_116,r77_117,r77_118,r77_119,r77_120,r77_121,r77_122,r77_123,r77_124,r77_125,r77_126,
	r78_0,r78_1,r78_2,r78_3,r78_4,r78_5,r78_6,r78_7,r78_8,r78_9,r78_10,r78_11,r78_12,r78_13,r78_14,r78_15,r78_16,
		r78_17,r78_18,r78_19,r78_20,r78_21,r78_22,r78_23,r78_24,r78_25,r78_26,r78_27,r78_28,r78_29,r78_30,r78_31,r78_32,
		r78_33,r78_34,r78_35,r78_36,r78_37,r78_38,r78_39,r78_40,r78_41,r78_42,r78_43,r78_44,r78_45,r78_46,r78_47,r78_48,
		r78_49,r78_50,r78_51,r78_52,r78_53,r78_54,r78_55,r78_56,r78_57,r78_58,r78_59,r78_60,r78_61,r78_62,r78_63,r78_64,
		r78_65,r78_66,r78_67,r78_68,r78_69,r78_70,r78_71,r78_72,r78_73,r78_74,r78_75,r78_76,r78_77,r78_78,r78_79,r78_80,
		r78_81,r78_82,r78_83,r78_84,r78_85,r78_86,r78_87,r78_88,r78_89,r78_90,r78_91,r78_92,r78_93,r78_94,r78_95,r78_96,
		r78_97,r78_98,r78_99,r78_100,r78_101,r78_102,r78_103,r78_104,r78_105,r78_106,r78_107,r78_108,r78_109,r78_110,r78_111,r78_112,
		r78_113,r78_114,r78_115,r78_116,r78_117,r78_118,r78_119,r78_120,r78_121,r78_122,r78_123,r78_124,r78_125,r78_126,
	r79_0,r79_1,r79_2,r79_3,r79_4,r79_5,r79_6,r79_7,r79_8,r79_9,r79_10,r79_11,r79_12,r79_13,r79_14,r79_15,r79_16,
		r79_17,r79_18,r79_19,r79_20,r79_21,r79_22,r79_23,r79_24,r79_25,r79_26,r79_27,r79_28,r79_29,r79_30,r79_31,r79_32,
		r79_33,r79_34,r79_35,r79_36,r79_37,r79_38,r79_39,r79_40,r79_41,r79_42,r79_43,r79_44,r79_45,r79_46,r79_47,r79_48,
		r79_49,r79_50,r79_51,r79_52,r79_53,r79_54,r79_55,r79_56,r79_57,r79_58,r79_59,r79_60,r79_61,r79_62,r79_63,r79_64,
		r79_65,r79_66,r79_67,r79_68,r79_69,r79_70,r79_71,r79_72,r79_73,r79_74,r79_75,r79_76,r79_77,r79_78,r79_79,r79_80,
		r79_81,r79_82,r79_83,r79_84,r79_85,r79_86,r79_87,r79_88,r79_89,r79_90,r79_91,r79_92,r79_93,r79_94,r79_95,r79_96,
		r79_97,r79_98,r79_99,r79_100,r79_101,r79_102,r79_103,r79_104,r79_105,r79_106,r79_107,r79_108,r79_109,r79_110,r79_111,r79_112,
		r79_113,r79_114,r79_115,r79_116,r79_117,r79_118,r79_119,r79_120,r79_121,r79_122,r79_123,r79_124,r79_125,r79_126,
	r80_0,r80_1,r80_2,r80_3,r80_4,r80_5,r80_6,r80_7,r80_8,r80_9,r80_10,r80_11,r80_12,r80_13,r80_14,r80_15,r80_16,
		r80_17,r80_18,r80_19,r80_20,r80_21,r80_22,r80_23,r80_24,r80_25,r80_26,r80_27,r80_28,r80_29,r80_30,r80_31,r80_32,
		r80_33,r80_34,r80_35,r80_36,r80_37,r80_38,r80_39,r80_40,r80_41,r80_42,r80_43,r80_44,r80_45,r80_46,r80_47,r80_48,
		r80_49,r80_50,r80_51,r80_52,r80_53,r80_54,r80_55,r80_56,r80_57,r80_58,r80_59,r80_60,r80_61,r80_62,r80_63,r80_64,
		r80_65,r80_66,r80_67,r80_68,r80_69,r80_70,r80_71,r80_72,r80_73,r80_74,r80_75,r80_76,r80_77,r80_78,r80_79,r80_80,
		r80_81,r80_82,r80_83,r80_84,r80_85,r80_86,r80_87,r80_88,r80_89,r80_90,r80_91,r80_92,r80_93,r80_94,r80_95,r80_96,
		r80_97,r80_98,r80_99,r80_100,r80_101,r80_102,r80_103,r80_104,r80_105,r80_106,r80_107,r80_108,r80_109,r80_110,r80_111,r80_112,
		r80_113,r80_114,r80_115,r80_116,r80_117,r80_118,r80_119,r80_120,r80_121,r80_122,r80_123,r80_124,r80_125,r80_126,
	r81_0,r81_1,r81_2,r81_3,r81_4,r81_5,r81_6,r81_7,r81_8,r81_9,r81_10,r81_11,r81_12,r81_13,r81_14,r81_15,r81_16,
		r81_17,r81_18,r81_19,r81_20,r81_21,r81_22,r81_23,r81_24,r81_25,r81_26,r81_27,r81_28,r81_29,r81_30,r81_31,r81_32,
		r81_33,r81_34,r81_35,r81_36,r81_37,r81_38,r81_39,r81_40,r81_41,r81_42,r81_43,r81_44,r81_45,r81_46,r81_47,r81_48,
		r81_49,r81_50,r81_51,r81_52,r81_53,r81_54,r81_55,r81_56,r81_57,r81_58,r81_59,r81_60,r81_61,r81_62,r81_63,r81_64,
		r81_65,r81_66,r81_67,r81_68,r81_69,r81_70,r81_71,r81_72,r81_73,r81_74,r81_75,r81_76,r81_77,r81_78,r81_79,r81_80,
		r81_81,r81_82,r81_83,r81_84,r81_85,r81_86,r81_87,r81_88,r81_89,r81_90,r81_91,r81_92,r81_93,r81_94,r81_95,r81_96,
		r81_97,r81_98,r81_99,r81_100,r81_101,r81_102,r81_103,r81_104,r81_105,r81_106,r81_107,r81_108,r81_109,r81_110,r81_111,r81_112,
		r81_113,r81_114,r81_115,r81_116,r81_117,r81_118,r81_119,r81_120,r81_121,r81_122,r81_123,r81_124,r81_125,r81_126,
	r82_0,r82_1,r82_2,r82_3,r82_4,r82_5,r82_6,r82_7,r82_8,r82_9,r82_10,r82_11,r82_12,r82_13,r82_14,r82_15,r82_16,
		r82_17,r82_18,r82_19,r82_20,r82_21,r82_22,r82_23,r82_24,r82_25,r82_26,r82_27,r82_28,r82_29,r82_30,r82_31,r82_32,
		r82_33,r82_34,r82_35,r82_36,r82_37,r82_38,r82_39,r82_40,r82_41,r82_42,r82_43,r82_44,r82_45,r82_46,r82_47,r82_48,
		r82_49,r82_50,r82_51,r82_52,r82_53,r82_54,r82_55,r82_56,r82_57,r82_58,r82_59,r82_60,r82_61,r82_62,r82_63,r82_64,
		r82_65,r82_66,r82_67,r82_68,r82_69,r82_70,r82_71,r82_72,r82_73,r82_74,r82_75,r82_76,r82_77,r82_78,r82_79,r82_80,
		r82_81,r82_82,r82_83,r82_84,r82_85,r82_86,r82_87,r82_88,r82_89,r82_90,r82_91,r82_92,r82_93,r82_94,r82_95,r82_96,
		r82_97,r82_98,r82_99,r82_100,r82_101,r82_102,r82_103,r82_104,r82_105,r82_106,r82_107,r82_108,r82_109,r82_110,r82_111,r82_112,
		r82_113,r82_114,r82_115,r82_116,r82_117,r82_118,r82_119,r82_120,r82_121,r82_122,r82_123,r82_124,r82_125,r82_126,
	r83_0,r83_1,r83_2,r83_3,r83_4,r83_5,r83_6,r83_7,r83_8,r83_9,r83_10,r83_11,r83_12,r83_13,r83_14,r83_15,r83_16,
		r83_17,r83_18,r83_19,r83_20,r83_21,r83_22,r83_23,r83_24,r83_25,r83_26,r83_27,r83_28,r83_29,r83_30,r83_31,r83_32,
		r83_33,r83_34,r83_35,r83_36,r83_37,r83_38,r83_39,r83_40,r83_41,r83_42,r83_43,r83_44,r83_45,r83_46,r83_47,r83_48,
		r83_49,r83_50,r83_51,r83_52,r83_53,r83_54,r83_55,r83_56,r83_57,r83_58,r83_59,r83_60,r83_61,r83_62,r83_63,r83_64,
		r83_65,r83_66,r83_67,r83_68,r83_69,r83_70,r83_71,r83_72,r83_73,r83_74,r83_75,r83_76,r83_77,r83_78,r83_79,r83_80,
		r83_81,r83_82,r83_83,r83_84,r83_85,r83_86,r83_87,r83_88,r83_89,r83_90,r83_91,r83_92,r83_93,r83_94,r83_95,r83_96,
		r83_97,r83_98,r83_99,r83_100,r83_101,r83_102,r83_103,r83_104,r83_105,r83_106,r83_107,r83_108,r83_109,r83_110,r83_111,r83_112,
		r83_113,r83_114,r83_115,r83_116,r83_117,r83_118,r83_119,r83_120,r83_121,r83_122,r83_123,r83_124,r83_125,r83_126,
	r84_0,r84_1,r84_2,r84_3,r84_4,r84_5,r84_6,r84_7,r84_8,r84_9,r84_10,r84_11,r84_12,r84_13,r84_14,r84_15,r84_16,
		r84_17,r84_18,r84_19,r84_20,r84_21,r84_22,r84_23,r84_24,r84_25,r84_26,r84_27,r84_28,r84_29,r84_30,r84_31,r84_32,
		r84_33,r84_34,r84_35,r84_36,r84_37,r84_38,r84_39,r84_40,r84_41,r84_42,r84_43,r84_44,r84_45,r84_46,r84_47,r84_48,
		r84_49,r84_50,r84_51,r84_52,r84_53,r84_54,r84_55,r84_56,r84_57,r84_58,r84_59,r84_60,r84_61,r84_62,r84_63,r84_64,
		r84_65,r84_66,r84_67,r84_68,r84_69,r84_70,r84_71,r84_72,r84_73,r84_74,r84_75,r84_76,r84_77,r84_78,r84_79,r84_80,
		r84_81,r84_82,r84_83,r84_84,r84_85,r84_86,r84_87,r84_88,r84_89,r84_90,r84_91,r84_92,r84_93,r84_94,r84_95,r84_96,
		r84_97,r84_98,r84_99,r84_100,r84_101,r84_102,r84_103,r84_104,r84_105,r84_106,r84_107,r84_108,r84_109,r84_110,r84_111,r84_112,
		r84_113,r84_114,r84_115,r84_116,r84_117,r84_118,r84_119,r84_120,r84_121,r84_122,r84_123,r84_124,r84_125,r84_126,
	r85_0,r85_1,r85_2,r85_3,r85_4,r85_5,r85_6,r85_7,r85_8,r85_9,r85_10,r85_11,r85_12,r85_13,r85_14,r85_15,r85_16,
		r85_17,r85_18,r85_19,r85_20,r85_21,r85_22,r85_23,r85_24,r85_25,r85_26,r85_27,r85_28,r85_29,r85_30,r85_31,r85_32,
		r85_33,r85_34,r85_35,r85_36,r85_37,r85_38,r85_39,r85_40,r85_41,r85_42,r85_43,r85_44,r85_45,r85_46,r85_47,r85_48,
		r85_49,r85_50,r85_51,r85_52,r85_53,r85_54,r85_55,r85_56,r85_57,r85_58,r85_59,r85_60,r85_61,r85_62,r85_63,r85_64,
		r85_65,r85_66,r85_67,r85_68,r85_69,r85_70,r85_71,r85_72,r85_73,r85_74,r85_75,r85_76,r85_77,r85_78,r85_79,r85_80,
		r85_81,r85_82,r85_83,r85_84,r85_85,r85_86,r85_87,r85_88,r85_89,r85_90,r85_91,r85_92,r85_93,r85_94,r85_95,r85_96,
		r85_97,r85_98,r85_99,r85_100,r85_101,r85_102,r85_103,r85_104,r85_105,r85_106,r85_107,r85_108,r85_109,r85_110,r85_111,r85_112,
		r85_113,r85_114,r85_115,r85_116,r85_117,r85_118,r85_119,r85_120,r85_121,r85_122,r85_123,r85_124,r85_125,r85_126,
	r86_0,r86_1,r86_2,r86_3,r86_4,r86_5,r86_6,r86_7,r86_8,r86_9,r86_10,r86_11,r86_12,r86_13,r86_14,r86_15,r86_16,
		r86_17,r86_18,r86_19,r86_20,r86_21,r86_22,r86_23,r86_24,r86_25,r86_26,r86_27,r86_28,r86_29,r86_30,r86_31,r86_32,
		r86_33,r86_34,r86_35,r86_36,r86_37,r86_38,r86_39,r86_40,r86_41,r86_42,r86_43,r86_44,r86_45,r86_46,r86_47,r86_48,
		r86_49,r86_50,r86_51,r86_52,r86_53,r86_54,r86_55,r86_56,r86_57,r86_58,r86_59,r86_60,r86_61,r86_62,r86_63,r86_64,
		r86_65,r86_66,r86_67,r86_68,r86_69,r86_70,r86_71,r86_72,r86_73,r86_74,r86_75,r86_76,r86_77,r86_78,r86_79,r86_80,
		r86_81,r86_82,r86_83,r86_84,r86_85,r86_86,r86_87,r86_88,r86_89,r86_90,r86_91,r86_92,r86_93,r86_94,r86_95,r86_96,
		r86_97,r86_98,r86_99,r86_100,r86_101,r86_102,r86_103,r86_104,r86_105,r86_106,r86_107,r86_108,r86_109,r86_110,r86_111,r86_112,
		r86_113,r86_114,r86_115,r86_116,r86_117,r86_118,r86_119,r86_120,r86_121,r86_122,r86_123,r86_124,r86_125,r86_126,
	r87_0,r87_1,r87_2,r87_3,r87_4,r87_5,r87_6,r87_7,r87_8,r87_9,r87_10,r87_11,r87_12,r87_13,r87_14,r87_15,r87_16,
		r87_17,r87_18,r87_19,r87_20,r87_21,r87_22,r87_23,r87_24,r87_25,r87_26,r87_27,r87_28,r87_29,r87_30,r87_31,r87_32,
		r87_33,r87_34,r87_35,r87_36,r87_37,r87_38,r87_39,r87_40,r87_41,r87_42,r87_43,r87_44,r87_45,r87_46,r87_47,r87_48,
		r87_49,r87_50,r87_51,r87_52,r87_53,r87_54,r87_55,r87_56,r87_57,r87_58,r87_59,r87_60,r87_61,r87_62,r87_63,r87_64,
		r87_65,r87_66,r87_67,r87_68,r87_69,r87_70,r87_71,r87_72,r87_73,r87_74,r87_75,r87_76,r87_77,r87_78,r87_79,r87_80,
		r87_81,r87_82,r87_83,r87_84,r87_85,r87_86,r87_87,r87_88,r87_89,r87_90,r87_91,r87_92,r87_93,r87_94,r87_95,r87_96,
		r87_97,r87_98,r87_99,r87_100,r87_101,r87_102,r87_103,r87_104,r87_105,r87_106,r87_107,r87_108,r87_109,r87_110,r87_111,r87_112,
		r87_113,r87_114,r87_115,r87_116,r87_117,r87_118,r87_119,r87_120,r87_121,r87_122,r87_123,r87_124,r87_125,r87_126,
	r88_0,r88_1,r88_2,r88_3,r88_4,r88_5,r88_6,r88_7,r88_8,r88_9,r88_10,r88_11,r88_12,r88_13,r88_14,r88_15,r88_16,
		r88_17,r88_18,r88_19,r88_20,r88_21,r88_22,r88_23,r88_24,r88_25,r88_26,r88_27,r88_28,r88_29,r88_30,r88_31,r88_32,
		r88_33,r88_34,r88_35,r88_36,r88_37,r88_38,r88_39,r88_40,r88_41,r88_42,r88_43,r88_44,r88_45,r88_46,r88_47,r88_48,
		r88_49,r88_50,r88_51,r88_52,r88_53,r88_54,r88_55,r88_56,r88_57,r88_58,r88_59,r88_60,r88_61,r88_62,r88_63,r88_64,
		r88_65,r88_66,r88_67,r88_68,r88_69,r88_70,r88_71,r88_72,r88_73,r88_74,r88_75,r88_76,r88_77,r88_78,r88_79,r88_80,
		r88_81,r88_82,r88_83,r88_84,r88_85,r88_86,r88_87,r88_88,r88_89,r88_90,r88_91,r88_92,r88_93,r88_94,r88_95,r88_96,
		r88_97,r88_98,r88_99,r88_100,r88_101,r88_102,r88_103,r88_104,r88_105,r88_106,r88_107,r88_108,r88_109,r88_110,r88_111,r88_112,
		r88_113,r88_114,r88_115,r88_116,r88_117,r88_118,r88_119,r88_120,r88_121,r88_122,r88_123,r88_124,r88_125,r88_126,
	r89_0,r89_1,r89_2,r89_3,r89_4,r89_5,r89_6,r89_7,r89_8,r89_9,r89_10,r89_11,r89_12,r89_13,r89_14,r89_15,r89_16,
		r89_17,r89_18,r89_19,r89_20,r89_21,r89_22,r89_23,r89_24,r89_25,r89_26,r89_27,r89_28,r89_29,r89_30,r89_31,r89_32,
		r89_33,r89_34,r89_35,r89_36,r89_37,r89_38,r89_39,r89_40,r89_41,r89_42,r89_43,r89_44,r89_45,r89_46,r89_47,r89_48,
		r89_49,r89_50,r89_51,r89_52,r89_53,r89_54,r89_55,r89_56,r89_57,r89_58,r89_59,r89_60,r89_61,r89_62,r89_63,r89_64,
		r89_65,r89_66,r89_67,r89_68,r89_69,r89_70,r89_71,r89_72,r89_73,r89_74,r89_75,r89_76,r89_77,r89_78,r89_79,r89_80,
		r89_81,r89_82,r89_83,r89_84,r89_85,r89_86,r89_87,r89_88,r89_89,r89_90,r89_91,r89_92,r89_93,r89_94,r89_95,r89_96,
		r89_97,r89_98,r89_99,r89_100,r89_101,r89_102,r89_103,r89_104,r89_105,r89_106,r89_107,r89_108,r89_109,r89_110,r89_111,r89_112,
		r89_113,r89_114,r89_115,r89_116,r89_117,r89_118,r89_119,r89_120,r89_121,r89_122,r89_123,r89_124,r89_125,r89_126,
	r90_0,r90_1,r90_2,r90_3,r90_4,r90_5,r90_6,r90_7,r90_8,r90_9,r90_10,r90_11,r90_12,r90_13,r90_14,r90_15,r90_16,
		r90_17,r90_18,r90_19,r90_20,r90_21,r90_22,r90_23,r90_24,r90_25,r90_26,r90_27,r90_28,r90_29,r90_30,r90_31,r90_32,
		r90_33,r90_34,r90_35,r90_36,r90_37,r90_38,r90_39,r90_40,r90_41,r90_42,r90_43,r90_44,r90_45,r90_46,r90_47,r90_48,
		r90_49,r90_50,r90_51,r90_52,r90_53,r90_54,r90_55,r90_56,r90_57,r90_58,r90_59,r90_60,r90_61,r90_62,r90_63,r90_64,
		r90_65,r90_66,r90_67,r90_68,r90_69,r90_70,r90_71,r90_72,r90_73,r90_74,r90_75,r90_76,r90_77,r90_78,r90_79,r90_80,
		r90_81,r90_82,r90_83,r90_84,r90_85,r90_86,r90_87,r90_88,r90_89,r90_90,r90_91,r90_92,r90_93,r90_94,r90_95,r90_96,
		r90_97,r90_98,r90_99,r90_100,r90_101,r90_102,r90_103,r90_104,r90_105,r90_106,r90_107,r90_108,r90_109,r90_110,r90_111,r90_112,
		r90_113,r90_114,r90_115,r90_116,r90_117,r90_118,r90_119,r90_120,r90_121,r90_122,r90_123,r90_124,r90_125,r90_126,
	r91_0,r91_1,r91_2,r91_3,r91_4,r91_5,r91_6,r91_7,r91_8,r91_9,r91_10,r91_11,r91_12,r91_13,r91_14,r91_15,r91_16,
		r91_17,r91_18,r91_19,r91_20,r91_21,r91_22,r91_23,r91_24,r91_25,r91_26,r91_27,r91_28,r91_29,r91_30,r91_31,r91_32,
		r91_33,r91_34,r91_35,r91_36,r91_37,r91_38,r91_39,r91_40,r91_41,r91_42,r91_43,r91_44,r91_45,r91_46,r91_47,r91_48,
		r91_49,r91_50,r91_51,r91_52,r91_53,r91_54,r91_55,r91_56,r91_57,r91_58,r91_59,r91_60,r91_61,r91_62,r91_63,r91_64,
		r91_65,r91_66,r91_67,r91_68,r91_69,r91_70,r91_71,r91_72,r91_73,r91_74,r91_75,r91_76,r91_77,r91_78,r91_79,r91_80,
		r91_81,r91_82,r91_83,r91_84,r91_85,r91_86,r91_87,r91_88,r91_89,r91_90,r91_91,r91_92,r91_93,r91_94,r91_95,r91_96,
		r91_97,r91_98,r91_99,r91_100,r91_101,r91_102,r91_103,r91_104,r91_105,r91_106,r91_107,r91_108,r91_109,r91_110,r91_111,r91_112,
		r91_113,r91_114,r91_115,r91_116,r91_117,r91_118,r91_119,r91_120,r91_121,r91_122,r91_123,r91_124,r91_125,r91_126,
	r92_0,r92_1,r92_2,r92_3,r92_4,r92_5,r92_6,r92_7,r92_8,r92_9,r92_10,r92_11,r92_12,r92_13,r92_14,r92_15,r92_16,
		r92_17,r92_18,r92_19,r92_20,r92_21,r92_22,r92_23,r92_24,r92_25,r92_26,r92_27,r92_28,r92_29,r92_30,r92_31,r92_32,
		r92_33,r92_34,r92_35,r92_36,r92_37,r92_38,r92_39,r92_40,r92_41,r92_42,r92_43,r92_44,r92_45,r92_46,r92_47,r92_48,
		r92_49,r92_50,r92_51,r92_52,r92_53,r92_54,r92_55,r92_56,r92_57,r92_58,r92_59,r92_60,r92_61,r92_62,r92_63,r92_64,
		r92_65,r92_66,r92_67,r92_68,r92_69,r92_70,r92_71,r92_72,r92_73,r92_74,r92_75,r92_76,r92_77,r92_78,r92_79,r92_80,
		r92_81,r92_82,r92_83,r92_84,r92_85,r92_86,r92_87,r92_88,r92_89,r92_90,r92_91,r92_92,r92_93,r92_94,r92_95,r92_96,
		r92_97,r92_98,r92_99,r92_100,r92_101,r92_102,r92_103,r92_104,r92_105,r92_106,r92_107,r92_108,r92_109,r92_110,r92_111,r92_112,
		r92_113,r92_114,r92_115,r92_116,r92_117,r92_118,r92_119,r92_120,r92_121,r92_122,r92_123,r92_124,r92_125,r92_126,
	r93_0,r93_1,r93_2,r93_3,r93_4,r93_5,r93_6,r93_7,r93_8,r93_9,r93_10,r93_11,r93_12,r93_13,r93_14,r93_15,r93_16,
		r93_17,r93_18,r93_19,r93_20,r93_21,r93_22,r93_23,r93_24,r93_25,r93_26,r93_27,r93_28,r93_29,r93_30,r93_31,r93_32,
		r93_33,r93_34,r93_35,r93_36,r93_37,r93_38,r93_39,r93_40,r93_41,r93_42,r93_43,r93_44,r93_45,r93_46,r93_47,r93_48,
		r93_49,r93_50,r93_51,r93_52,r93_53,r93_54,r93_55,r93_56,r93_57,r93_58,r93_59,r93_60,r93_61,r93_62,r93_63,r93_64,
		r93_65,r93_66,r93_67,r93_68,r93_69,r93_70,r93_71,r93_72,r93_73,r93_74,r93_75,r93_76,r93_77,r93_78,r93_79,r93_80,
		r93_81,r93_82,r93_83,r93_84,r93_85,r93_86,r93_87,r93_88,r93_89,r93_90,r93_91,r93_92,r93_93,r93_94,r93_95,r93_96,
		r93_97,r93_98,r93_99,r93_100,r93_101,r93_102,r93_103,r93_104,r93_105,r93_106,r93_107,r93_108,r93_109,r93_110,r93_111,r93_112,
		r93_113,r93_114,r93_115,r93_116,r93_117,r93_118,r93_119,r93_120,r93_121,r93_122,r93_123,r93_124,r93_125,r93_126,
	r94_0,r94_1,r94_2,r94_3,r94_4,r94_5,r94_6,r94_7,r94_8,r94_9,r94_10,r94_11,r94_12,r94_13,r94_14,r94_15,r94_16,
		r94_17,r94_18,r94_19,r94_20,r94_21,r94_22,r94_23,r94_24,r94_25,r94_26,r94_27,r94_28,r94_29,r94_30,r94_31,r94_32,
		r94_33,r94_34,r94_35,r94_36,r94_37,r94_38,r94_39,r94_40,r94_41,r94_42,r94_43,r94_44,r94_45,r94_46,r94_47,r94_48,
		r94_49,r94_50,r94_51,r94_52,r94_53,r94_54,r94_55,r94_56,r94_57,r94_58,r94_59,r94_60,r94_61,r94_62,r94_63,r94_64,
		r94_65,r94_66,r94_67,r94_68,r94_69,r94_70,r94_71,r94_72,r94_73,r94_74,r94_75,r94_76,r94_77,r94_78,r94_79,r94_80,
		r94_81,r94_82,r94_83,r94_84,r94_85,r94_86,r94_87,r94_88,r94_89,r94_90,r94_91,r94_92,r94_93,r94_94,r94_95,r94_96,
		r94_97,r94_98,r94_99,r94_100,r94_101,r94_102,r94_103,r94_104,r94_105,r94_106,r94_107,r94_108,r94_109,r94_110,r94_111,r94_112,
		r94_113,r94_114,r94_115,r94_116,r94_117,r94_118,r94_119,r94_120,r94_121,r94_122,r94_123,r94_124,r94_125,r94_126,
	r95_0,r95_1,r95_2,r95_3,r95_4,r95_5,r95_6,r95_7,r95_8,r95_9,r95_10,r95_11,r95_12,r95_13,r95_14,r95_15,r95_16,
		r95_17,r95_18,r95_19,r95_20,r95_21,r95_22,r95_23,r95_24,r95_25,r95_26,r95_27,r95_28,r95_29,r95_30,r95_31,r95_32,
		r95_33,r95_34,r95_35,r95_36,r95_37,r95_38,r95_39,r95_40,r95_41,r95_42,r95_43,r95_44,r95_45,r95_46,r95_47,r95_48,
		r95_49,r95_50,r95_51,r95_52,r95_53,r95_54,r95_55,r95_56,r95_57,r95_58,r95_59,r95_60,r95_61,r95_62,r95_63,r95_64,
		r95_65,r95_66,r95_67,r95_68,r95_69,r95_70,r95_71,r95_72,r95_73,r95_74,r95_75,r95_76,r95_77,r95_78,r95_79,r95_80,
		r95_81,r95_82,r95_83,r95_84,r95_85,r95_86,r95_87,r95_88,r95_89,r95_90,r95_91,r95_92,r95_93,r95_94,r95_95,r95_96,
		r95_97,r95_98,r95_99,r95_100,r95_101,r95_102,r95_103,r95_104,r95_105,r95_106,r95_107,r95_108,r95_109,r95_110,r95_111,r95_112,
		r95_113,r95_114,r95_115,r95_116,r95_117,r95_118,r95_119,r95_120,r95_121,r95_122,r95_123,r95_124,r95_125,r95_126,
	r96_0,r96_1,r96_2,r96_3,r96_4,r96_5,r96_6,r96_7,r96_8,r96_9,r96_10,r96_11,r96_12,r96_13,r96_14,r96_15,r96_16,
		r96_17,r96_18,r96_19,r96_20,r96_21,r96_22,r96_23,r96_24,r96_25,r96_26,r96_27,r96_28,r96_29,r96_30,r96_31,r96_32,
		r96_33,r96_34,r96_35,r96_36,r96_37,r96_38,r96_39,r96_40,r96_41,r96_42,r96_43,r96_44,r96_45,r96_46,r96_47,r96_48,
		r96_49,r96_50,r96_51,r96_52,r96_53,r96_54,r96_55,r96_56,r96_57,r96_58,r96_59,r96_60,r96_61,r96_62,r96_63,r96_64,
		r96_65,r96_66,r96_67,r96_68,r96_69,r96_70,r96_71,r96_72,r96_73,r96_74,r96_75,r96_76,r96_77,r96_78,r96_79,r96_80,
		r96_81,r96_82,r96_83,r96_84,r96_85,r96_86,r96_87,r96_88,r96_89,r96_90,r96_91,r96_92,r96_93,r96_94,r96_95,r96_96,
		r96_97,r96_98,r96_99,r96_100,r96_101,r96_102,r96_103,r96_104,r96_105,r96_106,r96_107,r96_108,r96_109,r96_110,r96_111,r96_112,
		r96_113,r96_114,r96_115,r96_116,r96_117,r96_118,r96_119,r96_120,r96_121,r96_122,r96_123,r96_124,r96_125,r96_126,
	r97_0,r97_1,r97_2,r97_3,r97_4,r97_5,r97_6,r97_7,r97_8,r97_9,r97_10,r97_11,r97_12,r97_13,r97_14,r97_15,r97_16,
		r97_17,r97_18,r97_19,r97_20,r97_21,r97_22,r97_23,r97_24,r97_25,r97_26,r97_27,r97_28,r97_29,r97_30,r97_31,r97_32,
		r97_33,r97_34,r97_35,r97_36,r97_37,r97_38,r97_39,r97_40,r97_41,r97_42,r97_43,r97_44,r97_45,r97_46,r97_47,r97_48,
		r97_49,r97_50,r97_51,r97_52,r97_53,r97_54,r97_55,r97_56,r97_57,r97_58,r97_59,r97_60,r97_61,r97_62,r97_63,r97_64,
		r97_65,r97_66,r97_67,r97_68,r97_69,r97_70,r97_71,r97_72,r97_73,r97_74,r97_75,r97_76,r97_77,r97_78,r97_79,r97_80,
		r97_81,r97_82,r97_83,r97_84,r97_85,r97_86,r97_87,r97_88,r97_89,r97_90,r97_91,r97_92,r97_93,r97_94,r97_95,r97_96,
		r97_97,r97_98,r97_99,r97_100,r97_101,r97_102,r97_103,r97_104,r97_105,r97_106,r97_107,r97_108,r97_109,r97_110,r97_111,r97_112,
		r97_113,r97_114,r97_115,r97_116,r97_117,r97_118,r97_119,r97_120,r97_121,r97_122,r97_123,r97_124,r97_125,r97_126,
	r98_0,r98_1,r98_2,r98_3,r98_4,r98_5,r98_6,r98_7,r98_8,r98_9,r98_10,r98_11,r98_12,r98_13,r98_14,r98_15,r98_16,
		r98_17,r98_18,r98_19,r98_20,r98_21,r98_22,r98_23,r98_24,r98_25,r98_26,r98_27,r98_28,r98_29,r98_30,r98_31,r98_32,
		r98_33,r98_34,r98_35,r98_36,r98_37,r98_38,r98_39,r98_40,r98_41,r98_42,r98_43,r98_44,r98_45,r98_46,r98_47,r98_48,
		r98_49,r98_50,r98_51,r98_52,r98_53,r98_54,r98_55,r98_56,r98_57,r98_58,r98_59,r98_60,r98_61,r98_62,r98_63,r98_64,
		r98_65,r98_66,r98_67,r98_68,r98_69,r98_70,r98_71,r98_72,r98_73,r98_74,r98_75,r98_76,r98_77,r98_78,r98_79,r98_80,
		r98_81,r98_82,r98_83,r98_84,r98_85,r98_86,r98_87,r98_88,r98_89,r98_90,r98_91,r98_92,r98_93,r98_94,r98_95,r98_96,
		r98_97,r98_98,r98_99,r98_100,r98_101,r98_102,r98_103,r98_104,r98_105,r98_106,r98_107,r98_108,r98_109,r98_110,r98_111,r98_112,
		r98_113,r98_114,r98_115,r98_116,r98_117,r98_118,r98_119,r98_120,r98_121,r98_122,r98_123,r98_124,r98_125,r98_126,
	r99_0,r99_1,r99_2,r99_3,r99_4,r99_5,r99_6,r99_7,r99_8,r99_9,r99_10,r99_11,r99_12,r99_13,r99_14,r99_15,r99_16,
		r99_17,r99_18,r99_19,r99_20,r99_21,r99_22,r99_23,r99_24,r99_25,r99_26,r99_27,r99_28,r99_29,r99_30,r99_31,r99_32,
		r99_33,r99_34,r99_35,r99_36,r99_37,r99_38,r99_39,r99_40,r99_41,r99_42,r99_43,r99_44,r99_45,r99_46,r99_47,r99_48,
		r99_49,r99_50,r99_51,r99_52,r99_53,r99_54,r99_55,r99_56,r99_57,r99_58,r99_59,r99_60,r99_61,r99_62,r99_63,r99_64,
		r99_65,r99_66,r99_67,r99_68,r99_69,r99_70,r99_71,r99_72,r99_73,r99_74,r99_75,r99_76,r99_77,r99_78,r99_79,r99_80,
		r99_81,r99_82,r99_83,r99_84,r99_85,r99_86,r99_87,r99_88,r99_89,r99_90,r99_91,r99_92,r99_93,r99_94,r99_95,r99_96,
		r99_97,r99_98,r99_99,r99_100,r99_101,r99_102,r99_103,r99_104,r99_105,r99_106,r99_107,r99_108,r99_109,r99_110,r99_111,r99_112,
		r99_113,r99_114,r99_115,r99_116,r99_117,r99_118,r99_119,r99_120,r99_121,r99_122,r99_123,r99_124,r99_125,r99_126,
	r100_0,r100_1,r100_2,r100_3,r100_4,r100_5,r100_6,r100_7,r100_8,r100_9,r100_10,r100_11,r100_12,r100_13,r100_14,r100_15,r100_16,
		r100_17,r100_18,r100_19,r100_20,r100_21,r100_22,r100_23,r100_24,r100_25,r100_26,r100_27,r100_28,r100_29,r100_30,r100_31,r100_32,
		r100_33,r100_34,r100_35,r100_36,r100_37,r100_38,r100_39,r100_40,r100_41,r100_42,r100_43,r100_44,r100_45,r100_46,r100_47,r100_48,
		r100_49,r100_50,r100_51,r100_52,r100_53,r100_54,r100_55,r100_56,r100_57,r100_58,r100_59,r100_60,r100_61,r100_62,r100_63,r100_64,
		r100_65,r100_66,r100_67,r100_68,r100_69,r100_70,r100_71,r100_72,r100_73,r100_74,r100_75,r100_76,r100_77,r100_78,r100_79,r100_80,
		r100_81,r100_82,r100_83,r100_84,r100_85,r100_86,r100_87,r100_88,r100_89,r100_90,r100_91,r100_92,r100_93,r100_94,r100_95,r100_96,
		r100_97,r100_98,r100_99,r100_100,r100_101,r100_102,r100_103,r100_104,r100_105,r100_106,r100_107,r100_108,r100_109,r100_110,r100_111,r100_112,
		r100_113,r100_114,r100_115,r100_116,r100_117,r100_118,r100_119,r100_120,r100_121,r100_122,r100_123,r100_124,r100_125,r100_126,
	r101_0,r101_1,r101_2,r101_3,r101_4,r101_5,r101_6,r101_7,r101_8,r101_9,r101_10,r101_11,r101_12,r101_13,r101_14,r101_15,r101_16,
		r101_17,r101_18,r101_19,r101_20,r101_21,r101_22,r101_23,r101_24,r101_25,r101_26,r101_27,r101_28,r101_29,r101_30,r101_31,r101_32,
		r101_33,r101_34,r101_35,r101_36,r101_37,r101_38,r101_39,r101_40,r101_41,r101_42,r101_43,r101_44,r101_45,r101_46,r101_47,r101_48,
		r101_49,r101_50,r101_51,r101_52,r101_53,r101_54,r101_55,r101_56,r101_57,r101_58,r101_59,r101_60,r101_61,r101_62,r101_63,r101_64,
		r101_65,r101_66,r101_67,r101_68,r101_69,r101_70,r101_71,r101_72,r101_73,r101_74,r101_75,r101_76,r101_77,r101_78,r101_79,r101_80,
		r101_81,r101_82,r101_83,r101_84,r101_85,r101_86,r101_87,r101_88,r101_89,r101_90,r101_91,r101_92,r101_93,r101_94,r101_95,r101_96,
		r101_97,r101_98,r101_99,r101_100,r101_101,r101_102,r101_103,r101_104,r101_105,r101_106,r101_107,r101_108,r101_109,r101_110,r101_111,r101_112,
		r101_113,r101_114,r101_115,r101_116,r101_117,r101_118,r101_119,r101_120,r101_121,r101_122,r101_123,r101_124,r101_125,r101_126,
	r102_0,r102_1,r102_2,r102_3,r102_4,r102_5,r102_6,r102_7,r102_8,r102_9,r102_10,r102_11,r102_12,r102_13,r102_14,r102_15,r102_16,
		r102_17,r102_18,r102_19,r102_20,r102_21,r102_22,r102_23,r102_24,r102_25,r102_26,r102_27,r102_28,r102_29,r102_30,r102_31,r102_32,
		r102_33,r102_34,r102_35,r102_36,r102_37,r102_38,r102_39,r102_40,r102_41,r102_42,r102_43,r102_44,r102_45,r102_46,r102_47,r102_48,
		r102_49,r102_50,r102_51,r102_52,r102_53,r102_54,r102_55,r102_56,r102_57,r102_58,r102_59,r102_60,r102_61,r102_62,r102_63,r102_64,
		r102_65,r102_66,r102_67,r102_68,r102_69,r102_70,r102_71,r102_72,r102_73,r102_74,r102_75,r102_76,r102_77,r102_78,r102_79,r102_80,
		r102_81,r102_82,r102_83,r102_84,r102_85,r102_86,r102_87,r102_88,r102_89,r102_90,r102_91,r102_92,r102_93,r102_94,r102_95,r102_96,
		r102_97,r102_98,r102_99,r102_100,r102_101,r102_102,r102_103,r102_104,r102_105,r102_106,r102_107,r102_108,r102_109,r102_110,r102_111,r102_112,
		r102_113,r102_114,r102_115,r102_116,r102_117,r102_118,r102_119,r102_120,r102_121,r102_122,r102_123,r102_124,r102_125,r102_126,
	r103_0,r103_1,r103_2,r103_3,r103_4,r103_5,r103_6,r103_7,r103_8,r103_9,r103_10,r103_11,r103_12,r103_13,r103_14,r103_15,r103_16,
		r103_17,r103_18,r103_19,r103_20,r103_21,r103_22,r103_23,r103_24,r103_25,r103_26,r103_27,r103_28,r103_29,r103_30,r103_31,r103_32,
		r103_33,r103_34,r103_35,r103_36,r103_37,r103_38,r103_39,r103_40,r103_41,r103_42,r103_43,r103_44,r103_45,r103_46,r103_47,r103_48,
		r103_49,r103_50,r103_51,r103_52,r103_53,r103_54,r103_55,r103_56,r103_57,r103_58,r103_59,r103_60,r103_61,r103_62,r103_63,r103_64,
		r103_65,r103_66,r103_67,r103_68,r103_69,r103_70,r103_71,r103_72,r103_73,r103_74,r103_75,r103_76,r103_77,r103_78,r103_79,r103_80,
		r103_81,r103_82,r103_83,r103_84,r103_85,r103_86,r103_87,r103_88,r103_89,r103_90,r103_91,r103_92,r103_93,r103_94,r103_95,r103_96,
		r103_97,r103_98,r103_99,r103_100,r103_101,r103_102,r103_103,r103_104,r103_105,r103_106,r103_107,r103_108,r103_109,r103_110,r103_111,r103_112,
		r103_113,r103_114,r103_115,r103_116,r103_117,r103_118,r103_119,r103_120,r103_121,r103_122,r103_123,r103_124,r103_125,r103_126,
	r104_0,r104_1,r104_2,r104_3,r104_4,r104_5,r104_6,r104_7,r104_8,r104_9,r104_10,r104_11,r104_12,r104_13,r104_14,r104_15,r104_16,
		r104_17,r104_18,r104_19,r104_20,r104_21,r104_22,r104_23,r104_24,r104_25,r104_26,r104_27,r104_28,r104_29,r104_30,r104_31,r104_32,
		r104_33,r104_34,r104_35,r104_36,r104_37,r104_38,r104_39,r104_40,r104_41,r104_42,r104_43,r104_44,r104_45,r104_46,r104_47,r104_48,
		r104_49,r104_50,r104_51,r104_52,r104_53,r104_54,r104_55,r104_56,r104_57,r104_58,r104_59,r104_60,r104_61,r104_62,r104_63,r104_64,
		r104_65,r104_66,r104_67,r104_68,r104_69,r104_70,r104_71,r104_72,r104_73,r104_74,r104_75,r104_76,r104_77,r104_78,r104_79,r104_80,
		r104_81,r104_82,r104_83,r104_84,r104_85,r104_86,r104_87,r104_88,r104_89,r104_90,r104_91,r104_92,r104_93,r104_94,r104_95,r104_96,
		r104_97,r104_98,r104_99,r104_100,r104_101,r104_102,r104_103,r104_104,r104_105,r104_106,r104_107,r104_108,r104_109,r104_110,r104_111,r104_112,
		r104_113,r104_114,r104_115,r104_116,r104_117,r104_118,r104_119,r104_120,r104_121,r104_122,r104_123,r104_124,r104_125,r104_126,
	r105_0,r105_1,r105_2,r105_3,r105_4,r105_5,r105_6,r105_7,r105_8,r105_9,r105_10,r105_11,r105_12,r105_13,r105_14,r105_15,r105_16,
		r105_17,r105_18,r105_19,r105_20,r105_21,r105_22,r105_23,r105_24,r105_25,r105_26,r105_27,r105_28,r105_29,r105_30,r105_31,r105_32,
		r105_33,r105_34,r105_35,r105_36,r105_37,r105_38,r105_39,r105_40,r105_41,r105_42,r105_43,r105_44,r105_45,r105_46,r105_47,r105_48,
		r105_49,r105_50,r105_51,r105_52,r105_53,r105_54,r105_55,r105_56,r105_57,r105_58,r105_59,r105_60,r105_61,r105_62,r105_63,r105_64,
		r105_65,r105_66,r105_67,r105_68,r105_69,r105_70,r105_71,r105_72,r105_73,r105_74,r105_75,r105_76,r105_77,r105_78,r105_79,r105_80,
		r105_81,r105_82,r105_83,r105_84,r105_85,r105_86,r105_87,r105_88,r105_89,r105_90,r105_91,r105_92,r105_93,r105_94,r105_95,r105_96,
		r105_97,r105_98,r105_99,r105_100,r105_101,r105_102,r105_103,r105_104,r105_105,r105_106,r105_107,r105_108,r105_109,r105_110,r105_111,r105_112,
		r105_113,r105_114,r105_115,r105_116,r105_117,r105_118,r105_119,r105_120,r105_121,r105_122,r105_123,r105_124,r105_125,r105_126,
	r106_0,r106_1,r106_2,r106_3,r106_4,r106_5,r106_6,r106_7,r106_8,r106_9,r106_10,r106_11,r106_12,r106_13,r106_14,r106_15,r106_16,
		r106_17,r106_18,r106_19,r106_20,r106_21,r106_22,r106_23,r106_24,r106_25,r106_26,r106_27,r106_28,r106_29,r106_30,r106_31,r106_32,
		r106_33,r106_34,r106_35,r106_36,r106_37,r106_38,r106_39,r106_40,r106_41,r106_42,r106_43,r106_44,r106_45,r106_46,r106_47,r106_48,
		r106_49,r106_50,r106_51,r106_52,r106_53,r106_54,r106_55,r106_56,r106_57,r106_58,r106_59,r106_60,r106_61,r106_62,r106_63,r106_64,
		r106_65,r106_66,r106_67,r106_68,r106_69,r106_70,r106_71,r106_72,r106_73,r106_74,r106_75,r106_76,r106_77,r106_78,r106_79,r106_80,
		r106_81,r106_82,r106_83,r106_84,r106_85,r106_86,r106_87,r106_88,r106_89,r106_90,r106_91,r106_92,r106_93,r106_94,r106_95,r106_96,
		r106_97,r106_98,r106_99,r106_100,r106_101,r106_102,r106_103,r106_104,r106_105,r106_106,r106_107,r106_108,r106_109,r106_110,r106_111,r106_112,
		r106_113,r106_114,r106_115,r106_116,r106_117,r106_118,r106_119,r106_120,r106_121,r106_122,r106_123,r106_124,r106_125,r106_126,
	r107_0,r107_1,r107_2,r107_3,r107_4,r107_5,r107_6,r107_7,r107_8,r107_9,r107_10,r107_11,r107_12,r107_13,r107_14,r107_15,r107_16,
		r107_17,r107_18,r107_19,r107_20,r107_21,r107_22,r107_23,r107_24,r107_25,r107_26,r107_27,r107_28,r107_29,r107_30,r107_31,r107_32,
		r107_33,r107_34,r107_35,r107_36,r107_37,r107_38,r107_39,r107_40,r107_41,r107_42,r107_43,r107_44,r107_45,r107_46,r107_47,r107_48,
		r107_49,r107_50,r107_51,r107_52,r107_53,r107_54,r107_55,r107_56,r107_57,r107_58,r107_59,r107_60,r107_61,r107_62,r107_63,r107_64,
		r107_65,r107_66,r107_67,r107_68,r107_69,r107_70,r107_71,r107_72,r107_73,r107_74,r107_75,r107_76,r107_77,r107_78,r107_79,r107_80,
		r107_81,r107_82,r107_83,r107_84,r107_85,r107_86,r107_87,r107_88,r107_89,r107_90,r107_91,r107_92,r107_93,r107_94,r107_95,r107_96,
		r107_97,r107_98,r107_99,r107_100,r107_101,r107_102,r107_103,r107_104,r107_105,r107_106,r107_107,r107_108,r107_109,r107_110,r107_111,r107_112,
		r107_113,r107_114,r107_115,r107_116,r107_117,r107_118,r107_119,r107_120,r107_121,r107_122,r107_123,r107_124,r107_125,r107_126,
	r108_0,r108_1,r108_2,r108_3,r108_4,r108_5,r108_6,r108_7,r108_8,r108_9,r108_10,r108_11,r108_12,r108_13,r108_14,r108_15,r108_16,
		r108_17,r108_18,r108_19,r108_20,r108_21,r108_22,r108_23,r108_24,r108_25,r108_26,r108_27,r108_28,r108_29,r108_30,r108_31,r108_32,
		r108_33,r108_34,r108_35,r108_36,r108_37,r108_38,r108_39,r108_40,r108_41,r108_42,r108_43,r108_44,r108_45,r108_46,r108_47,r108_48,
		r108_49,r108_50,r108_51,r108_52,r108_53,r108_54,r108_55,r108_56,r108_57,r108_58,r108_59,r108_60,r108_61,r108_62,r108_63,r108_64,
		r108_65,r108_66,r108_67,r108_68,r108_69,r108_70,r108_71,r108_72,r108_73,r108_74,r108_75,r108_76,r108_77,r108_78,r108_79,r108_80,
		r108_81,r108_82,r108_83,r108_84,r108_85,r108_86,r108_87,r108_88,r108_89,r108_90,r108_91,r108_92,r108_93,r108_94,r108_95,r108_96,
		r108_97,r108_98,r108_99,r108_100,r108_101,r108_102,r108_103,r108_104,r108_105,r108_106,r108_107,r108_108,r108_109,r108_110,r108_111,r108_112,
		r108_113,r108_114,r108_115,r108_116,r108_117,r108_118,r108_119,r108_120,r108_121,r108_122,r108_123,r108_124,r108_125,r108_126,
	r109_0,r109_1,r109_2,r109_3,r109_4,r109_5,r109_6,r109_7,r109_8,r109_9,r109_10,r109_11,r109_12,r109_13,r109_14,r109_15,r109_16,
		r109_17,r109_18,r109_19,r109_20,r109_21,r109_22,r109_23,r109_24,r109_25,r109_26,r109_27,r109_28,r109_29,r109_30,r109_31,r109_32,
		r109_33,r109_34,r109_35,r109_36,r109_37,r109_38,r109_39,r109_40,r109_41,r109_42,r109_43,r109_44,r109_45,r109_46,r109_47,r109_48,
		r109_49,r109_50,r109_51,r109_52,r109_53,r109_54,r109_55,r109_56,r109_57,r109_58,r109_59,r109_60,r109_61,r109_62,r109_63,r109_64,
		r109_65,r109_66,r109_67,r109_68,r109_69,r109_70,r109_71,r109_72,r109_73,r109_74,r109_75,r109_76,r109_77,r109_78,r109_79,r109_80,
		r109_81,r109_82,r109_83,r109_84,r109_85,r109_86,r109_87,r109_88,r109_89,r109_90,r109_91,r109_92,r109_93,r109_94,r109_95,r109_96,
		r109_97,r109_98,r109_99,r109_100,r109_101,r109_102,r109_103,r109_104,r109_105,r109_106,r109_107,r109_108,r109_109,r109_110,r109_111,r109_112,
		r109_113,r109_114,r109_115,r109_116,r109_117,r109_118,r109_119,r109_120,r109_121,r109_122,r109_123,r109_124,r109_125,r109_126,
	r110_0,r110_1,r110_2,r110_3,r110_4,r110_5,r110_6,r110_7,r110_8,r110_9,r110_10,r110_11,r110_12,r110_13,r110_14,r110_15,r110_16,
		r110_17,r110_18,r110_19,r110_20,r110_21,r110_22,r110_23,r110_24,r110_25,r110_26,r110_27,r110_28,r110_29,r110_30,r110_31,r110_32,
		r110_33,r110_34,r110_35,r110_36,r110_37,r110_38,r110_39,r110_40,r110_41,r110_42,r110_43,r110_44,r110_45,r110_46,r110_47,r110_48,
		r110_49,r110_50,r110_51,r110_52,r110_53,r110_54,r110_55,r110_56,r110_57,r110_58,r110_59,r110_60,r110_61,r110_62,r110_63,r110_64,
		r110_65,r110_66,r110_67,r110_68,r110_69,r110_70,r110_71,r110_72,r110_73,r110_74,r110_75,r110_76,r110_77,r110_78,r110_79,r110_80,
		r110_81,r110_82,r110_83,r110_84,r110_85,r110_86,r110_87,r110_88,r110_89,r110_90,r110_91,r110_92,r110_93,r110_94,r110_95,r110_96,
		r110_97,r110_98,r110_99,r110_100,r110_101,r110_102,r110_103,r110_104,r110_105,r110_106,r110_107,r110_108,r110_109,r110_110,r110_111,r110_112,
		r110_113,r110_114,r110_115,r110_116,r110_117,r110_118,r110_119,r110_120,r110_121,r110_122,r110_123,r110_124,r110_125,r110_126,
	r111_0,r111_1,r111_2,r111_3,r111_4,r111_5,r111_6,r111_7,r111_8,r111_9,r111_10,r111_11,r111_12,r111_13,r111_14,r111_15,r111_16,
		r111_17,r111_18,r111_19,r111_20,r111_21,r111_22,r111_23,r111_24,r111_25,r111_26,r111_27,r111_28,r111_29,r111_30,r111_31,r111_32,
		r111_33,r111_34,r111_35,r111_36,r111_37,r111_38,r111_39,r111_40,r111_41,r111_42,r111_43,r111_44,r111_45,r111_46,r111_47,r111_48,
		r111_49,r111_50,r111_51,r111_52,r111_53,r111_54,r111_55,r111_56,r111_57,r111_58,r111_59,r111_60,r111_61,r111_62,r111_63,r111_64,
		r111_65,r111_66,r111_67,r111_68,r111_69,r111_70,r111_71,r111_72,r111_73,r111_74,r111_75,r111_76,r111_77,r111_78,r111_79,r111_80,
		r111_81,r111_82,r111_83,r111_84,r111_85,r111_86,r111_87,r111_88,r111_89,r111_90,r111_91,r111_92,r111_93,r111_94,r111_95,r111_96,
		r111_97,r111_98,r111_99,r111_100,r111_101,r111_102,r111_103,r111_104,r111_105,r111_106,r111_107,r111_108,r111_109,r111_110,r111_111,r111_112,
		r111_113,r111_114,r111_115,r111_116,r111_117,r111_118,r111_119,r111_120,r111_121,r111_122,r111_123,r111_124,r111_125,r111_126,
	r112_0,r112_1,r112_2,r112_3,r112_4,r112_5,r112_6,r112_7,r112_8,r112_9,r112_10,r112_11,r112_12,r112_13,r112_14,r112_15,r112_16,
		r112_17,r112_18,r112_19,r112_20,r112_21,r112_22,r112_23,r112_24,r112_25,r112_26,r112_27,r112_28,r112_29,r112_30,r112_31,r112_32,
		r112_33,r112_34,r112_35,r112_36,r112_37,r112_38,r112_39,r112_40,r112_41,r112_42,r112_43,r112_44,r112_45,r112_46,r112_47,r112_48,
		r112_49,r112_50,r112_51,r112_52,r112_53,r112_54,r112_55,r112_56,r112_57,r112_58,r112_59,r112_60,r112_61,r112_62,r112_63,r112_64,
		r112_65,r112_66,r112_67,r112_68,r112_69,r112_70,r112_71,r112_72,r112_73,r112_74,r112_75,r112_76,r112_77,r112_78,r112_79,r112_80,
		r112_81,r112_82,r112_83,r112_84,r112_85,r112_86,r112_87,r112_88,r112_89,r112_90,r112_91,r112_92,r112_93,r112_94,r112_95,r112_96,
		r112_97,r112_98,r112_99,r112_100,r112_101,r112_102,r112_103,r112_104,r112_105,r112_106,r112_107,r112_108,r112_109,r112_110,r112_111,r112_112,
		r112_113,r112_114,r112_115,r112_116,r112_117,r112_118,r112_119,r112_120,r112_121,r112_122,r112_123,r112_124,r112_125,r112_126,
	r113_0,r113_1,r113_2,r113_3,r113_4,r113_5,r113_6,r113_7,r113_8,r113_9,r113_10,r113_11,r113_12,r113_13,r113_14,r113_15,r113_16,
		r113_17,r113_18,r113_19,r113_20,r113_21,r113_22,r113_23,r113_24,r113_25,r113_26,r113_27,r113_28,r113_29,r113_30,r113_31,r113_32,
		r113_33,r113_34,r113_35,r113_36,r113_37,r113_38,r113_39,r113_40,r113_41,r113_42,r113_43,r113_44,r113_45,r113_46,r113_47,r113_48,
		r113_49,r113_50,r113_51,r113_52,r113_53,r113_54,r113_55,r113_56,r113_57,r113_58,r113_59,r113_60,r113_61,r113_62,r113_63,r113_64,
		r113_65,r113_66,r113_67,r113_68,r113_69,r113_70,r113_71,r113_72,r113_73,r113_74,r113_75,r113_76,r113_77,r113_78,r113_79,r113_80,
		r113_81,r113_82,r113_83,r113_84,r113_85,r113_86,r113_87,r113_88,r113_89,r113_90,r113_91,r113_92,r113_93,r113_94,r113_95,r113_96,
		r113_97,r113_98,r113_99,r113_100,r113_101,r113_102,r113_103,r113_104,r113_105,r113_106,r113_107,r113_108,r113_109,r113_110,r113_111,r113_112,
		r113_113,r113_114,r113_115,r113_116,r113_117,r113_118,r113_119,r113_120,r113_121,r113_122,r113_123,r113_124,r113_125,r113_126,
	r114_0,r114_1,r114_2,r114_3,r114_4,r114_5,r114_6,r114_7,r114_8,r114_9,r114_10,r114_11,r114_12,r114_13,r114_14,r114_15,r114_16,
		r114_17,r114_18,r114_19,r114_20,r114_21,r114_22,r114_23,r114_24,r114_25,r114_26,r114_27,r114_28,r114_29,r114_30,r114_31,r114_32,
		r114_33,r114_34,r114_35,r114_36,r114_37,r114_38,r114_39,r114_40,r114_41,r114_42,r114_43,r114_44,r114_45,r114_46,r114_47,r114_48,
		r114_49,r114_50,r114_51,r114_52,r114_53,r114_54,r114_55,r114_56,r114_57,r114_58,r114_59,r114_60,r114_61,r114_62,r114_63,r114_64,
		r114_65,r114_66,r114_67,r114_68,r114_69,r114_70,r114_71,r114_72,r114_73,r114_74,r114_75,r114_76,r114_77,r114_78,r114_79,r114_80,
		r114_81,r114_82,r114_83,r114_84,r114_85,r114_86,r114_87,r114_88,r114_89,r114_90,r114_91,r114_92,r114_93,r114_94,r114_95,r114_96,
		r114_97,r114_98,r114_99,r114_100,r114_101,r114_102,r114_103,r114_104,r114_105,r114_106,r114_107,r114_108,r114_109,r114_110,r114_111,r114_112,
		r114_113,r114_114,r114_115,r114_116,r114_117,r114_118,r114_119,r114_120,r114_121,r114_122,r114_123,r114_124,r114_125,r114_126,
	r115_0,r115_1,r115_2,r115_3,r115_4,r115_5,r115_6,r115_7,r115_8,r115_9,r115_10,r115_11,r115_12,r115_13,r115_14,r115_15,r115_16,
		r115_17,r115_18,r115_19,r115_20,r115_21,r115_22,r115_23,r115_24,r115_25,r115_26,r115_27,r115_28,r115_29,r115_30,r115_31,r115_32,
		r115_33,r115_34,r115_35,r115_36,r115_37,r115_38,r115_39,r115_40,r115_41,r115_42,r115_43,r115_44,r115_45,r115_46,r115_47,r115_48,
		r115_49,r115_50,r115_51,r115_52,r115_53,r115_54,r115_55,r115_56,r115_57,r115_58,r115_59,r115_60,r115_61,r115_62,r115_63,r115_64,
		r115_65,r115_66,r115_67,r115_68,r115_69,r115_70,r115_71,r115_72,r115_73,r115_74,r115_75,r115_76,r115_77,r115_78,r115_79,r115_80,
		r115_81,r115_82,r115_83,r115_84,r115_85,r115_86,r115_87,r115_88,r115_89,r115_90,r115_91,r115_92,r115_93,r115_94,r115_95,r115_96,
		r115_97,r115_98,r115_99,r115_100,r115_101,r115_102,r115_103,r115_104,r115_105,r115_106,r115_107,r115_108,r115_109,r115_110,r115_111,r115_112,
		r115_113,r115_114,r115_115,r115_116,r115_117,r115_118,r115_119,r115_120,r115_121,r115_122,r115_123,r115_124,r115_125,r115_126,
	r116_0,r116_1,r116_2,r116_3,r116_4,r116_5,r116_6,r116_7,r116_8,r116_9,r116_10,r116_11,r116_12,r116_13,r116_14,r116_15,r116_16,
		r116_17,r116_18,r116_19,r116_20,r116_21,r116_22,r116_23,r116_24,r116_25,r116_26,r116_27,r116_28,r116_29,r116_30,r116_31,r116_32,
		r116_33,r116_34,r116_35,r116_36,r116_37,r116_38,r116_39,r116_40,r116_41,r116_42,r116_43,r116_44,r116_45,r116_46,r116_47,r116_48,
		r116_49,r116_50,r116_51,r116_52,r116_53,r116_54,r116_55,r116_56,r116_57,r116_58,r116_59,r116_60,r116_61,r116_62,r116_63,r116_64,
		r116_65,r116_66,r116_67,r116_68,r116_69,r116_70,r116_71,r116_72,r116_73,r116_74,r116_75,r116_76,r116_77,r116_78,r116_79,r116_80,
		r116_81,r116_82,r116_83,r116_84,r116_85,r116_86,r116_87,r116_88,r116_89,r116_90,r116_91,r116_92,r116_93,r116_94,r116_95,r116_96,
		r116_97,r116_98,r116_99,r116_100,r116_101,r116_102,r116_103,r116_104,r116_105,r116_106,r116_107,r116_108,r116_109,r116_110,r116_111,r116_112,
		r116_113,r116_114,r116_115,r116_116,r116_117,r116_118,r116_119,r116_120,r116_121,r116_122,r116_123,r116_124,r116_125,r116_126,
	r117_0,r117_1,r117_2,r117_3,r117_4,r117_5,r117_6,r117_7,r117_8,r117_9,r117_10,r117_11,r117_12,r117_13,r117_14,r117_15,r117_16,
		r117_17,r117_18,r117_19,r117_20,r117_21,r117_22,r117_23,r117_24,r117_25,r117_26,r117_27,r117_28,r117_29,r117_30,r117_31,r117_32,
		r117_33,r117_34,r117_35,r117_36,r117_37,r117_38,r117_39,r117_40,r117_41,r117_42,r117_43,r117_44,r117_45,r117_46,r117_47,r117_48,
		r117_49,r117_50,r117_51,r117_52,r117_53,r117_54,r117_55,r117_56,r117_57,r117_58,r117_59,r117_60,r117_61,r117_62,r117_63,r117_64,
		r117_65,r117_66,r117_67,r117_68,r117_69,r117_70,r117_71,r117_72,r117_73,r117_74,r117_75,r117_76,r117_77,r117_78,r117_79,r117_80,
		r117_81,r117_82,r117_83,r117_84,r117_85,r117_86,r117_87,r117_88,r117_89,r117_90,r117_91,r117_92,r117_93,r117_94,r117_95,r117_96,
		r117_97,r117_98,r117_99,r117_100,r117_101,r117_102,r117_103,r117_104,r117_105,r117_106,r117_107,r117_108,r117_109,r117_110,r117_111,r117_112,
		r117_113,r117_114,r117_115,r117_116,r117_117,r117_118,r117_119,r117_120,r117_121,r117_122,r117_123,r117_124,r117_125,r117_126,
	r118_0,r118_1,r118_2,r118_3,r118_4,r118_5,r118_6,r118_7,r118_8,r118_9,r118_10,r118_11,r118_12,r118_13,r118_14,r118_15,r118_16,
		r118_17,r118_18,r118_19,r118_20,r118_21,r118_22,r118_23,r118_24,r118_25,r118_26,r118_27,r118_28,r118_29,r118_30,r118_31,r118_32,
		r118_33,r118_34,r118_35,r118_36,r118_37,r118_38,r118_39,r118_40,r118_41,r118_42,r118_43,r118_44,r118_45,r118_46,r118_47,r118_48,
		r118_49,r118_50,r118_51,r118_52,r118_53,r118_54,r118_55,r118_56,r118_57,r118_58,r118_59,r118_60,r118_61,r118_62,r118_63,r118_64,
		r118_65,r118_66,r118_67,r118_68,r118_69,r118_70,r118_71,r118_72,r118_73,r118_74,r118_75,r118_76,r118_77,r118_78,r118_79,r118_80,
		r118_81,r118_82,r118_83,r118_84,r118_85,r118_86,r118_87,r118_88,r118_89,r118_90,r118_91,r118_92,r118_93,r118_94,r118_95,r118_96,
		r118_97,r118_98,r118_99,r118_100,r118_101,r118_102,r118_103,r118_104,r118_105,r118_106,r118_107,r118_108,r118_109,r118_110,r118_111,r118_112,
		r118_113,r118_114,r118_115,r118_116,r118_117,r118_118,r118_119,r118_120,r118_121,r118_122,r118_123,r118_124,r118_125,r118_126,
	r119_0,r119_1,r119_2,r119_3,r119_4,r119_5,r119_6,r119_7,r119_8,r119_9,r119_10,r119_11,r119_12,r119_13,r119_14,r119_15,r119_16,
		r119_17,r119_18,r119_19,r119_20,r119_21,r119_22,r119_23,r119_24,r119_25,r119_26,r119_27,r119_28,r119_29,r119_30,r119_31,r119_32,
		r119_33,r119_34,r119_35,r119_36,r119_37,r119_38,r119_39,r119_40,r119_41,r119_42,r119_43,r119_44,r119_45,r119_46,r119_47,r119_48,
		r119_49,r119_50,r119_51,r119_52,r119_53,r119_54,r119_55,r119_56,r119_57,r119_58,r119_59,r119_60,r119_61,r119_62,r119_63,r119_64,
		r119_65,r119_66,r119_67,r119_68,r119_69,r119_70,r119_71,r119_72,r119_73,r119_74,r119_75,r119_76,r119_77,r119_78,r119_79,r119_80,
		r119_81,r119_82,r119_83,r119_84,r119_85,r119_86,r119_87,r119_88,r119_89,r119_90,r119_91,r119_92,r119_93,r119_94,r119_95,r119_96,
		r119_97,r119_98,r119_99,r119_100,r119_101,r119_102,r119_103,r119_104,r119_105,r119_106,r119_107,r119_108,r119_109,r119_110,r119_111,r119_112,
		r119_113,r119_114,r119_115,r119_116,r119_117,r119_118,r119_119,r119_120,r119_121,r119_122,r119_123,r119_124,r119_125,r119_126,
	r120_0,r120_1,r120_2,r120_3,r120_4,r120_5,r120_6,r120_7,r120_8,r120_9,r120_10,r120_11,r120_12,r120_13,r120_14,r120_15,r120_16,
		r120_17,r120_18,r120_19,r120_20,r120_21,r120_22,r120_23,r120_24,r120_25,r120_26,r120_27,r120_28,r120_29,r120_30,r120_31,r120_32,
		r120_33,r120_34,r120_35,r120_36,r120_37,r120_38,r120_39,r120_40,r120_41,r120_42,r120_43,r120_44,r120_45,r120_46,r120_47,r120_48,
		r120_49,r120_50,r120_51,r120_52,r120_53,r120_54,r120_55,r120_56,r120_57,r120_58,r120_59,r120_60,r120_61,r120_62,r120_63,r120_64,
		r120_65,r120_66,r120_67,r120_68,r120_69,r120_70,r120_71,r120_72,r120_73,r120_74,r120_75,r120_76,r120_77,r120_78,r120_79,r120_80,
		r120_81,r120_82,r120_83,r120_84,r120_85,r120_86,r120_87,r120_88,r120_89,r120_90,r120_91,r120_92,r120_93,r120_94,r120_95,r120_96,
		r120_97,r120_98,r120_99,r120_100,r120_101,r120_102,r120_103,r120_104,r120_105,r120_106,r120_107,r120_108,r120_109,r120_110,r120_111,r120_112,
		r120_113,r120_114,r120_115,r120_116,r120_117,r120_118,r120_119,r120_120,r120_121,r120_122,r120_123,r120_124,r120_125,r120_126,
	r121_0,r121_1,r121_2,r121_3,r121_4,r121_5,r121_6,r121_7,r121_8,r121_9,r121_10,r121_11,r121_12,r121_13,r121_14,r121_15,r121_16,
		r121_17,r121_18,r121_19,r121_20,r121_21,r121_22,r121_23,r121_24,r121_25,r121_26,r121_27,r121_28,r121_29,r121_30,r121_31,r121_32,
		r121_33,r121_34,r121_35,r121_36,r121_37,r121_38,r121_39,r121_40,r121_41,r121_42,r121_43,r121_44,r121_45,r121_46,r121_47,r121_48,
		r121_49,r121_50,r121_51,r121_52,r121_53,r121_54,r121_55,r121_56,r121_57,r121_58,r121_59,r121_60,r121_61,r121_62,r121_63,r121_64,
		r121_65,r121_66,r121_67,r121_68,r121_69,r121_70,r121_71,r121_72,r121_73,r121_74,r121_75,r121_76,r121_77,r121_78,r121_79,r121_80,
		r121_81,r121_82,r121_83,r121_84,r121_85,r121_86,r121_87,r121_88,r121_89,r121_90,r121_91,r121_92,r121_93,r121_94,r121_95,r121_96,
		r121_97,r121_98,r121_99,r121_100,r121_101,r121_102,r121_103,r121_104,r121_105,r121_106,r121_107,r121_108,r121_109,r121_110,r121_111,r121_112,
		r121_113,r121_114,r121_115,r121_116,r121_117,r121_118,r121_119,r121_120,r121_121,r121_122,r121_123,r121_124,r121_125,r121_126,
	r122_0,r122_1,r122_2,r122_3,r122_4,r122_5,r122_6,r122_7,r122_8,r122_9,r122_10,r122_11,r122_12,r122_13,r122_14,r122_15,r122_16,
		r122_17,r122_18,r122_19,r122_20,r122_21,r122_22,r122_23,r122_24,r122_25,r122_26,r122_27,r122_28,r122_29,r122_30,r122_31,r122_32,
		r122_33,r122_34,r122_35,r122_36,r122_37,r122_38,r122_39,r122_40,r122_41,r122_42,r122_43,r122_44,r122_45,r122_46,r122_47,r122_48,
		r122_49,r122_50,r122_51,r122_52,r122_53,r122_54,r122_55,r122_56,r122_57,r122_58,r122_59,r122_60,r122_61,r122_62,r122_63,r122_64,
		r122_65,r122_66,r122_67,r122_68,r122_69,r122_70,r122_71,r122_72,r122_73,r122_74,r122_75,r122_76,r122_77,r122_78,r122_79,r122_80,
		r122_81,r122_82,r122_83,r122_84,r122_85,r122_86,r122_87,r122_88,r122_89,r122_90,r122_91,r122_92,r122_93,r122_94,r122_95,r122_96,
		r122_97,r122_98,r122_99,r122_100,r122_101,r122_102,r122_103,r122_104,r122_105,r122_106,r122_107,r122_108,r122_109,r122_110,r122_111,r122_112,
		r122_113,r122_114,r122_115,r122_116,r122_117,r122_118,r122_119,r122_120,r122_121,r122_122,r122_123,r122_124,r122_125,r122_126,
	r123_0,r123_1,r123_2,r123_3,r123_4,r123_5,r123_6,r123_7,r123_8,r123_9,r123_10,r123_11,r123_12,r123_13,r123_14,r123_15,r123_16,
		r123_17,r123_18,r123_19,r123_20,r123_21,r123_22,r123_23,r123_24,r123_25,r123_26,r123_27,r123_28,r123_29,r123_30,r123_31,r123_32,
		r123_33,r123_34,r123_35,r123_36,r123_37,r123_38,r123_39,r123_40,r123_41,r123_42,r123_43,r123_44,r123_45,r123_46,r123_47,r123_48,
		r123_49,r123_50,r123_51,r123_52,r123_53,r123_54,r123_55,r123_56,r123_57,r123_58,r123_59,r123_60,r123_61,r123_62,r123_63,r123_64,
		r123_65,r123_66,r123_67,r123_68,r123_69,r123_70,r123_71,r123_72,r123_73,r123_74,r123_75,r123_76,r123_77,r123_78,r123_79,r123_80,
		r123_81,r123_82,r123_83,r123_84,r123_85,r123_86,r123_87,r123_88,r123_89,r123_90,r123_91,r123_92,r123_93,r123_94,r123_95,r123_96,
		r123_97,r123_98,r123_99,r123_100,r123_101,r123_102,r123_103,r123_104,r123_105,r123_106,r123_107,r123_108,r123_109,r123_110,r123_111,r123_112,
		r123_113,r123_114,r123_115,r123_116,r123_117,r123_118,r123_119,r123_120,r123_121,r123_122,r123_123,r123_124,r123_125,r123_126,
	r124_0,r124_1,r124_2,r124_3,r124_4,r124_5,r124_6,r124_7,r124_8,r124_9,r124_10,r124_11,r124_12,r124_13,r124_14,r124_15,r124_16,
		r124_17,r124_18,r124_19,r124_20,r124_21,r124_22,r124_23,r124_24,r124_25,r124_26,r124_27,r124_28,r124_29,r124_30,r124_31,r124_32,
		r124_33,r124_34,r124_35,r124_36,r124_37,r124_38,r124_39,r124_40,r124_41,r124_42,r124_43,r124_44,r124_45,r124_46,r124_47,r124_48,
		r124_49,r124_50,r124_51,r124_52,r124_53,r124_54,r124_55,r124_56,r124_57,r124_58,r124_59,r124_60,r124_61,r124_62,r124_63,r124_64,
		r124_65,r124_66,r124_67,r124_68,r124_69,r124_70,r124_71,r124_72,r124_73,r124_74,r124_75,r124_76,r124_77,r124_78,r124_79,r124_80,
		r124_81,r124_82,r124_83,r124_84,r124_85,r124_86,r124_87,r124_88,r124_89,r124_90,r124_91,r124_92,r124_93,r124_94,r124_95,r124_96,
		r124_97,r124_98,r124_99,r124_100,r124_101,r124_102,r124_103,r124_104,r124_105,r124_106,r124_107,r124_108,r124_109,r124_110,r124_111,r124_112,
		r124_113,r124_114,r124_115,r124_116,r124_117,r124_118,r124_119,r124_120,r124_121,r124_122,r124_123,r124_124,r124_125,r124_126,
	r125_0,r125_1,r125_2,r125_3,r125_4,r125_5,r125_6,r125_7,r125_8,r125_9,r125_10,r125_11,r125_12,r125_13,r125_14,r125_15,r125_16,
		r125_17,r125_18,r125_19,r125_20,r125_21,r125_22,r125_23,r125_24,r125_25,r125_26,r125_27,r125_28,r125_29,r125_30,r125_31,r125_32,
		r125_33,r125_34,r125_35,r125_36,r125_37,r125_38,r125_39,r125_40,r125_41,r125_42,r125_43,r125_44,r125_45,r125_46,r125_47,r125_48,
		r125_49,r125_50,r125_51,r125_52,r125_53,r125_54,r125_55,r125_56,r125_57,r125_58,r125_59,r125_60,r125_61,r125_62,r125_63,r125_64,
		r125_65,r125_66,r125_67,r125_68,r125_69,r125_70,r125_71,r125_72,r125_73,r125_74,r125_75,r125_76,r125_77,r125_78,r125_79,r125_80,
		r125_81,r125_82,r125_83,r125_84,r125_85,r125_86,r125_87,r125_88,r125_89,r125_90,r125_91,r125_92,r125_93,r125_94,r125_95,r125_96,
		r125_97,r125_98,r125_99,r125_100,r125_101,r125_102,r125_103,r125_104,r125_105,r125_106,r125_107,r125_108,r125_109,r125_110,r125_111,r125_112,
		r125_113,r125_114,r125_115,r125_116,r125_117,r125_118,r125_119,r125_120,r125_121,r125_122,r125_123,r125_124,r125_125,r125_126,
	r126_0,r126_1,r126_2,r126_3,r126_4,r126_5,r126_6,r126_7,r126_8,r126_9,r126_10,r126_11,r126_12,r126_13,r126_14,r126_15,r126_16,
		r126_17,r126_18,r126_19,r126_20,r126_21,r126_22,r126_23,r126_24,r126_25,r126_26,r126_27,r126_28,r126_29,r126_30,r126_31,r126_32,
		r126_33,r126_34,r126_35,r126_36,r126_37,r126_38,r126_39,r126_40,r126_41,r126_42,r126_43,r126_44,r126_45,r126_46,r126_47,r126_48,
		r126_49,r126_50,r126_51,r126_52,r126_53,r126_54,r126_55,r126_56,r126_57,r126_58,r126_59,r126_60,r126_61,r126_62,r126_63,r126_64,
		r126_65,r126_66,r126_67,r126_68,r126_69,r126_70,r126_71,r126_72,r126_73,r126_74,r126_75,r126_76,r126_77,r126_78,r126_79,r126_80,
		r126_81,r126_82,r126_83,r126_84,r126_85,r126_86,r126_87,r126_88,r126_89,r126_90,r126_91,r126_92,r126_93,r126_94,r126_95,r126_96,
		r126_97,r126_98,r126_99,r126_100,r126_101,r126_102,r126_103,r126_104,r126_105,r126_106,r126_107,r126_108,r126_109,r126_110,r126_111,r126_112,
		r126_113,r126_114,r126_115,r126_116,r126_117,r126_118,r126_119,r126_120,r126_121,r126_122,r126_123,r126_124,r126_125,r126_126,
	r127_0,r127_1,r127_2,r127_3,r127_4,r127_5,r127_6,r127_7,r127_8,r127_9,r127_10,r127_11,r127_12,r127_13,r127_14,r127_15,r127_16,
		r127_17,r127_18,r127_19,r127_20,r127_21,r127_22,r127_23,r127_24,r127_25,r127_26,r127_27,r127_28,r127_29,r127_30,r127_31,r127_32,
		r127_33,r127_34,r127_35,r127_36,r127_37,r127_38,r127_39,r127_40,r127_41,r127_42,r127_43,r127_44,r127_45,r127_46,r127_47,r127_48,
		r127_49,r127_50,r127_51,r127_52,r127_53,r127_54,r127_55,r127_56,r127_57,r127_58,r127_59,r127_60,r127_61,r127_62,r127_63,r127_64,
		r127_65,r127_66,r127_67,r127_68,r127_69,r127_70,r127_71,r127_72,r127_73,r127_74,r127_75,r127_76,r127_77,r127_78,r127_79,r127_80,
		r127_81,r127_82,r127_83,r127_84,r127_85,r127_86,r127_87,r127_88,r127_89,r127_90,r127_91,r127_92,r127_93,r127_94,r127_95,r127_96,
		r127_97,r127_98,r127_99,r127_100,r127_101,r127_102,r127_103,r127_104,r127_105,r127_106,r127_107,r127_108,r127_109,r127_110,r127_111,r127_112,
		r127_113,r127_114,r127_115,r127_116,r127_117,r127_118,r127_119,r127_120,r127_121,r127_122,r127_123,r127_124,r127_125,r127_126;
	

	PE pe0_0(.x(x0),.w(w0),.acc(32'h0),.res(r0_0),.clk(clk),.wout(w0_0));
	PE pe0_1(.x(x1),.w(w0_0),.acc(r0_0),.res(r0_1),.clk(clk),.wout(w0_1));
	PE pe0_2(.x(x2),.w(w0_1),.acc(r0_1),.res(r0_2),.clk(clk),.wout(w0_2));
	PE pe0_3(.x(x3),.w(w0_2),.acc(r0_2),.res(r0_3),.clk(clk),.wout(w0_3));
	PE pe0_4(.x(x4),.w(w0_3),.acc(r0_3),.res(r0_4),.clk(clk),.wout(w0_4));
	PE pe0_5(.x(x5),.w(w0_4),.acc(r0_4),.res(r0_5),.clk(clk),.wout(w0_5));
	PE pe0_6(.x(x6),.w(w0_5),.acc(r0_5),.res(r0_6),.clk(clk),.wout(w0_6));
	PE pe0_7(.x(x7),.w(w0_6),.acc(r0_6),.res(r0_7),.clk(clk),.wout(w0_7));
	PE pe0_8(.x(x8),.w(w0_7),.acc(r0_7),.res(r0_8),.clk(clk),.wout(w0_8));
	PE pe0_9(.x(x9),.w(w0_8),.acc(r0_8),.res(r0_9),.clk(clk),.wout(w0_9));
	PE pe0_10(.x(x10),.w(w0_9),.acc(r0_9),.res(r0_10),.clk(clk),.wout(w0_10));
	PE pe0_11(.x(x11),.w(w0_10),.acc(r0_10),.res(r0_11),.clk(clk),.wout(w0_11));
	PE pe0_12(.x(x12),.w(w0_11),.acc(r0_11),.res(r0_12),.clk(clk),.wout(w0_12));
	PE pe0_13(.x(x13),.w(w0_12),.acc(r0_12),.res(r0_13),.clk(clk),.wout(w0_13));
	PE pe0_14(.x(x14),.w(w0_13),.acc(r0_13),.res(r0_14),.clk(clk),.wout(w0_14));
	PE pe0_15(.x(x15),.w(w0_14),.acc(r0_14),.res(r0_15),.clk(clk),.wout(w0_15));
	PE pe0_16(.x(x16),.w(w0_15),.acc(r0_15),.res(r0_16),.clk(clk),.wout(w0_16));
	PE pe0_17(.x(x17),.w(w0_16),.acc(r0_16),.res(r0_17),.clk(clk),.wout(w0_17));
	PE pe0_18(.x(x18),.w(w0_17),.acc(r0_17),.res(r0_18),.clk(clk),.wout(w0_18));
	PE pe0_19(.x(x19),.w(w0_18),.acc(r0_18),.res(r0_19),.clk(clk),.wout(w0_19));
	PE pe0_20(.x(x20),.w(w0_19),.acc(r0_19),.res(r0_20),.clk(clk),.wout(w0_20));
	PE pe0_21(.x(x21),.w(w0_20),.acc(r0_20),.res(r0_21),.clk(clk),.wout(w0_21));
	PE pe0_22(.x(x22),.w(w0_21),.acc(r0_21),.res(r0_22),.clk(clk),.wout(w0_22));
	PE pe0_23(.x(x23),.w(w0_22),.acc(r0_22),.res(r0_23),.clk(clk),.wout(w0_23));
	PE pe0_24(.x(x24),.w(w0_23),.acc(r0_23),.res(r0_24),.clk(clk),.wout(w0_24));
	PE pe0_25(.x(x25),.w(w0_24),.acc(r0_24),.res(r0_25),.clk(clk),.wout(w0_25));
	PE pe0_26(.x(x26),.w(w0_25),.acc(r0_25),.res(r0_26),.clk(clk),.wout(w0_26));
	PE pe0_27(.x(x27),.w(w0_26),.acc(r0_26),.res(r0_27),.clk(clk),.wout(w0_27));
	PE pe0_28(.x(x28),.w(w0_27),.acc(r0_27),.res(r0_28),.clk(clk),.wout(w0_28));
	PE pe0_29(.x(x29),.w(w0_28),.acc(r0_28),.res(r0_29),.clk(clk),.wout(w0_29));
	PE pe0_30(.x(x30),.w(w0_29),.acc(r0_29),.res(r0_30),.clk(clk),.wout(w0_30));
	PE pe0_31(.x(x31),.w(w0_30),.acc(r0_30),.res(r0_31),.clk(clk),.wout(w0_31));
	PE pe0_32(.x(x32),.w(w0_31),.acc(r0_31),.res(r0_32),.clk(clk),.wout(w0_32));
	PE pe0_33(.x(x33),.w(w0_32),.acc(r0_32),.res(r0_33),.clk(clk),.wout(w0_33));
	PE pe0_34(.x(x34),.w(w0_33),.acc(r0_33),.res(r0_34),.clk(clk),.wout(w0_34));
	PE pe0_35(.x(x35),.w(w0_34),.acc(r0_34),.res(r0_35),.clk(clk),.wout(w0_35));
	PE pe0_36(.x(x36),.w(w0_35),.acc(r0_35),.res(r0_36),.clk(clk),.wout(w0_36));
	PE pe0_37(.x(x37),.w(w0_36),.acc(r0_36),.res(r0_37),.clk(clk),.wout(w0_37));
	PE pe0_38(.x(x38),.w(w0_37),.acc(r0_37),.res(r0_38),.clk(clk),.wout(w0_38));
	PE pe0_39(.x(x39),.w(w0_38),.acc(r0_38),.res(r0_39),.clk(clk),.wout(w0_39));
	PE pe0_40(.x(x40),.w(w0_39),.acc(r0_39),.res(r0_40),.clk(clk),.wout(w0_40));
	PE pe0_41(.x(x41),.w(w0_40),.acc(r0_40),.res(r0_41),.clk(clk),.wout(w0_41));
	PE pe0_42(.x(x42),.w(w0_41),.acc(r0_41),.res(r0_42),.clk(clk),.wout(w0_42));
	PE pe0_43(.x(x43),.w(w0_42),.acc(r0_42),.res(r0_43),.clk(clk),.wout(w0_43));
	PE pe0_44(.x(x44),.w(w0_43),.acc(r0_43),.res(r0_44),.clk(clk),.wout(w0_44));
	PE pe0_45(.x(x45),.w(w0_44),.acc(r0_44),.res(r0_45),.clk(clk),.wout(w0_45));
	PE pe0_46(.x(x46),.w(w0_45),.acc(r0_45),.res(r0_46),.clk(clk),.wout(w0_46));
	PE pe0_47(.x(x47),.w(w0_46),.acc(r0_46),.res(r0_47),.clk(clk),.wout(w0_47));
	PE pe0_48(.x(x48),.w(w0_47),.acc(r0_47),.res(r0_48),.clk(clk),.wout(w0_48));
	PE pe0_49(.x(x49),.w(w0_48),.acc(r0_48),.res(r0_49),.clk(clk),.wout(w0_49));
	PE pe0_50(.x(x50),.w(w0_49),.acc(r0_49),.res(r0_50),.clk(clk),.wout(w0_50));
	PE pe0_51(.x(x51),.w(w0_50),.acc(r0_50),.res(r0_51),.clk(clk),.wout(w0_51));
	PE pe0_52(.x(x52),.w(w0_51),.acc(r0_51),.res(r0_52),.clk(clk),.wout(w0_52));
	PE pe0_53(.x(x53),.w(w0_52),.acc(r0_52),.res(r0_53),.clk(clk),.wout(w0_53));
	PE pe0_54(.x(x54),.w(w0_53),.acc(r0_53),.res(r0_54),.clk(clk),.wout(w0_54));
	PE pe0_55(.x(x55),.w(w0_54),.acc(r0_54),.res(r0_55),.clk(clk),.wout(w0_55));
	PE pe0_56(.x(x56),.w(w0_55),.acc(r0_55),.res(r0_56),.clk(clk),.wout(w0_56));
	PE pe0_57(.x(x57),.w(w0_56),.acc(r0_56),.res(r0_57),.clk(clk),.wout(w0_57));
	PE pe0_58(.x(x58),.w(w0_57),.acc(r0_57),.res(r0_58),.clk(clk),.wout(w0_58));
	PE pe0_59(.x(x59),.w(w0_58),.acc(r0_58),.res(r0_59),.clk(clk),.wout(w0_59));
	PE pe0_60(.x(x60),.w(w0_59),.acc(r0_59),.res(r0_60),.clk(clk),.wout(w0_60));
	PE pe0_61(.x(x61),.w(w0_60),.acc(r0_60),.res(r0_61),.clk(clk),.wout(w0_61));
	PE pe0_62(.x(x62),.w(w0_61),.acc(r0_61),.res(r0_62),.clk(clk),.wout(w0_62));
	PE pe0_63(.x(x63),.w(w0_62),.acc(r0_62),.res(r0_63),.clk(clk),.wout(w0_63));
	PE pe0_64(.x(x64),.w(w0_63),.acc(r0_63),.res(r0_64),.clk(clk),.wout(w0_64));
	PE pe0_65(.x(x65),.w(w0_64),.acc(r0_64),.res(r0_65),.clk(clk),.wout(w0_65));
	PE pe0_66(.x(x66),.w(w0_65),.acc(r0_65),.res(r0_66),.clk(clk),.wout(w0_66));
	PE pe0_67(.x(x67),.w(w0_66),.acc(r0_66),.res(r0_67),.clk(clk),.wout(w0_67));
	PE pe0_68(.x(x68),.w(w0_67),.acc(r0_67),.res(r0_68),.clk(clk),.wout(w0_68));
	PE pe0_69(.x(x69),.w(w0_68),.acc(r0_68),.res(r0_69),.clk(clk),.wout(w0_69));
	PE pe0_70(.x(x70),.w(w0_69),.acc(r0_69),.res(r0_70),.clk(clk),.wout(w0_70));
	PE pe0_71(.x(x71),.w(w0_70),.acc(r0_70),.res(r0_71),.clk(clk),.wout(w0_71));
	PE pe0_72(.x(x72),.w(w0_71),.acc(r0_71),.res(r0_72),.clk(clk),.wout(w0_72));
	PE pe0_73(.x(x73),.w(w0_72),.acc(r0_72),.res(r0_73),.clk(clk),.wout(w0_73));
	PE pe0_74(.x(x74),.w(w0_73),.acc(r0_73),.res(r0_74),.clk(clk),.wout(w0_74));
	PE pe0_75(.x(x75),.w(w0_74),.acc(r0_74),.res(r0_75),.clk(clk),.wout(w0_75));
	PE pe0_76(.x(x76),.w(w0_75),.acc(r0_75),.res(r0_76),.clk(clk),.wout(w0_76));
	PE pe0_77(.x(x77),.w(w0_76),.acc(r0_76),.res(r0_77),.clk(clk),.wout(w0_77));
	PE pe0_78(.x(x78),.w(w0_77),.acc(r0_77),.res(r0_78),.clk(clk),.wout(w0_78));
	PE pe0_79(.x(x79),.w(w0_78),.acc(r0_78),.res(r0_79),.clk(clk),.wout(w0_79));
	PE pe0_80(.x(x80),.w(w0_79),.acc(r0_79),.res(r0_80),.clk(clk),.wout(w0_80));
	PE pe0_81(.x(x81),.w(w0_80),.acc(r0_80),.res(r0_81),.clk(clk),.wout(w0_81));
	PE pe0_82(.x(x82),.w(w0_81),.acc(r0_81),.res(r0_82),.clk(clk),.wout(w0_82));
	PE pe0_83(.x(x83),.w(w0_82),.acc(r0_82),.res(r0_83),.clk(clk),.wout(w0_83));
	PE pe0_84(.x(x84),.w(w0_83),.acc(r0_83),.res(r0_84),.clk(clk),.wout(w0_84));
	PE pe0_85(.x(x85),.w(w0_84),.acc(r0_84),.res(r0_85),.clk(clk),.wout(w0_85));
	PE pe0_86(.x(x86),.w(w0_85),.acc(r0_85),.res(r0_86),.clk(clk),.wout(w0_86));
	PE pe0_87(.x(x87),.w(w0_86),.acc(r0_86),.res(r0_87),.clk(clk),.wout(w0_87));
	PE pe0_88(.x(x88),.w(w0_87),.acc(r0_87),.res(r0_88),.clk(clk),.wout(w0_88));
	PE pe0_89(.x(x89),.w(w0_88),.acc(r0_88),.res(r0_89),.clk(clk),.wout(w0_89));
	PE pe0_90(.x(x90),.w(w0_89),.acc(r0_89),.res(r0_90),.clk(clk),.wout(w0_90));
	PE pe0_91(.x(x91),.w(w0_90),.acc(r0_90),.res(r0_91),.clk(clk),.wout(w0_91));
	PE pe0_92(.x(x92),.w(w0_91),.acc(r0_91),.res(r0_92),.clk(clk),.wout(w0_92));
	PE pe0_93(.x(x93),.w(w0_92),.acc(r0_92),.res(r0_93),.clk(clk),.wout(w0_93));
	PE pe0_94(.x(x94),.w(w0_93),.acc(r0_93),.res(r0_94),.clk(clk),.wout(w0_94));
	PE pe0_95(.x(x95),.w(w0_94),.acc(r0_94),.res(r0_95),.clk(clk),.wout(w0_95));
	PE pe0_96(.x(x96),.w(w0_95),.acc(r0_95),.res(r0_96),.clk(clk),.wout(w0_96));
	PE pe0_97(.x(x97),.w(w0_96),.acc(r0_96),.res(r0_97),.clk(clk),.wout(w0_97));
	PE pe0_98(.x(x98),.w(w0_97),.acc(r0_97),.res(r0_98),.clk(clk),.wout(w0_98));
	PE pe0_99(.x(x99),.w(w0_98),.acc(r0_98),.res(r0_99),.clk(clk),.wout(w0_99));
	PE pe0_100(.x(x100),.w(w0_99),.acc(r0_99),.res(r0_100),.clk(clk),.wout(w0_100));
	PE pe0_101(.x(x101),.w(w0_100),.acc(r0_100),.res(r0_101),.clk(clk),.wout(w0_101));
	PE pe0_102(.x(x102),.w(w0_101),.acc(r0_101),.res(r0_102),.clk(clk),.wout(w0_102));
	PE pe0_103(.x(x103),.w(w0_102),.acc(r0_102),.res(r0_103),.clk(clk),.wout(w0_103));
	PE pe0_104(.x(x104),.w(w0_103),.acc(r0_103),.res(r0_104),.clk(clk),.wout(w0_104));
	PE pe0_105(.x(x105),.w(w0_104),.acc(r0_104),.res(r0_105),.clk(clk),.wout(w0_105));
	PE pe0_106(.x(x106),.w(w0_105),.acc(r0_105),.res(r0_106),.clk(clk),.wout(w0_106));
	PE pe0_107(.x(x107),.w(w0_106),.acc(r0_106),.res(r0_107),.clk(clk),.wout(w0_107));
	PE pe0_108(.x(x108),.w(w0_107),.acc(r0_107),.res(r0_108),.clk(clk),.wout(w0_108));
	PE pe0_109(.x(x109),.w(w0_108),.acc(r0_108),.res(r0_109),.clk(clk),.wout(w0_109));
	PE pe0_110(.x(x110),.w(w0_109),.acc(r0_109),.res(r0_110),.clk(clk),.wout(w0_110));
	PE pe0_111(.x(x111),.w(w0_110),.acc(r0_110),.res(r0_111),.clk(clk),.wout(w0_111));
	PE pe0_112(.x(x112),.w(w0_111),.acc(r0_111),.res(r0_112),.clk(clk),.wout(w0_112));
	PE pe0_113(.x(x113),.w(w0_112),.acc(r0_112),.res(r0_113),.clk(clk),.wout(w0_113));
	PE pe0_114(.x(x114),.w(w0_113),.acc(r0_113),.res(r0_114),.clk(clk),.wout(w0_114));
	PE pe0_115(.x(x115),.w(w0_114),.acc(r0_114),.res(r0_115),.clk(clk),.wout(w0_115));
	PE pe0_116(.x(x116),.w(w0_115),.acc(r0_115),.res(r0_116),.clk(clk),.wout(w0_116));
	PE pe0_117(.x(x117),.w(w0_116),.acc(r0_116),.res(r0_117),.clk(clk),.wout(w0_117));
	PE pe0_118(.x(x118),.w(w0_117),.acc(r0_117),.res(r0_118),.clk(clk),.wout(w0_118));
	PE pe0_119(.x(x119),.w(w0_118),.acc(r0_118),.res(r0_119),.clk(clk),.wout(w0_119));
	PE pe0_120(.x(x120),.w(w0_119),.acc(r0_119),.res(r0_120),.clk(clk),.wout(w0_120));
	PE pe0_121(.x(x121),.w(w0_120),.acc(r0_120),.res(r0_121),.clk(clk),.wout(w0_121));
	PE pe0_122(.x(x122),.w(w0_121),.acc(r0_121),.res(r0_122),.clk(clk),.wout(w0_122));
	PE pe0_123(.x(x123),.w(w0_122),.acc(r0_122),.res(r0_123),.clk(clk),.wout(w0_123));
	PE pe0_124(.x(x124),.w(w0_123),.acc(r0_123),.res(r0_124),.clk(clk),.wout(w0_124));
	PE pe0_125(.x(x125),.w(w0_124),.acc(r0_124),.res(r0_125),.clk(clk),.wout(w0_125));
	PE pe0_126(.x(x126),.w(w0_125),.acc(r0_125),.res(r0_126),.clk(clk),.wout(w0_126));
	PE pe0_127(.x(x127),.w(w0_126),.acc(r0_126),.res(result0),.clk(clk),.wout(weight0));

	PE pe1_0(.x(x0),.w(w1),.acc(32'h0),.res(r1_0),.clk(clk),.wout(w1_0));
	PE pe1_1(.x(x1),.w(w1_0),.acc(r1_0),.res(r1_1),.clk(clk),.wout(w1_1));
	PE pe1_2(.x(x2),.w(w1_1),.acc(r1_1),.res(r1_2),.clk(clk),.wout(w1_2));
	PE pe1_3(.x(x3),.w(w1_2),.acc(r1_2),.res(r1_3),.clk(clk),.wout(w1_3));
	PE pe1_4(.x(x4),.w(w1_3),.acc(r1_3),.res(r1_4),.clk(clk),.wout(w1_4));
	PE pe1_5(.x(x5),.w(w1_4),.acc(r1_4),.res(r1_5),.clk(clk),.wout(w1_5));
	PE pe1_6(.x(x6),.w(w1_5),.acc(r1_5),.res(r1_6),.clk(clk),.wout(w1_6));
	PE pe1_7(.x(x7),.w(w1_6),.acc(r1_6),.res(r1_7),.clk(clk),.wout(w1_7));
	PE pe1_8(.x(x8),.w(w1_7),.acc(r1_7),.res(r1_8),.clk(clk),.wout(w1_8));
	PE pe1_9(.x(x9),.w(w1_8),.acc(r1_8),.res(r1_9),.clk(clk),.wout(w1_9));
	PE pe1_10(.x(x10),.w(w1_9),.acc(r1_9),.res(r1_10),.clk(clk),.wout(w1_10));
	PE pe1_11(.x(x11),.w(w1_10),.acc(r1_10),.res(r1_11),.clk(clk),.wout(w1_11));
	PE pe1_12(.x(x12),.w(w1_11),.acc(r1_11),.res(r1_12),.clk(clk),.wout(w1_12));
	PE pe1_13(.x(x13),.w(w1_12),.acc(r1_12),.res(r1_13),.clk(clk),.wout(w1_13));
	PE pe1_14(.x(x14),.w(w1_13),.acc(r1_13),.res(r1_14),.clk(clk),.wout(w1_14));
	PE pe1_15(.x(x15),.w(w1_14),.acc(r1_14),.res(r1_15),.clk(clk),.wout(w1_15));
	PE pe1_16(.x(x16),.w(w1_15),.acc(r1_15),.res(r1_16),.clk(clk),.wout(w1_16));
	PE pe1_17(.x(x17),.w(w1_16),.acc(r1_16),.res(r1_17),.clk(clk),.wout(w1_17));
	PE pe1_18(.x(x18),.w(w1_17),.acc(r1_17),.res(r1_18),.clk(clk),.wout(w1_18));
	PE pe1_19(.x(x19),.w(w1_18),.acc(r1_18),.res(r1_19),.clk(clk),.wout(w1_19));
	PE pe1_20(.x(x20),.w(w1_19),.acc(r1_19),.res(r1_20),.clk(clk),.wout(w1_20));
	PE pe1_21(.x(x21),.w(w1_20),.acc(r1_20),.res(r1_21),.clk(clk),.wout(w1_21));
	PE pe1_22(.x(x22),.w(w1_21),.acc(r1_21),.res(r1_22),.clk(clk),.wout(w1_22));
	PE pe1_23(.x(x23),.w(w1_22),.acc(r1_22),.res(r1_23),.clk(clk),.wout(w1_23));
	PE pe1_24(.x(x24),.w(w1_23),.acc(r1_23),.res(r1_24),.clk(clk),.wout(w1_24));
	PE pe1_25(.x(x25),.w(w1_24),.acc(r1_24),.res(r1_25),.clk(clk),.wout(w1_25));
	PE pe1_26(.x(x26),.w(w1_25),.acc(r1_25),.res(r1_26),.clk(clk),.wout(w1_26));
	PE pe1_27(.x(x27),.w(w1_26),.acc(r1_26),.res(r1_27),.clk(clk),.wout(w1_27));
	PE pe1_28(.x(x28),.w(w1_27),.acc(r1_27),.res(r1_28),.clk(clk),.wout(w1_28));
	PE pe1_29(.x(x29),.w(w1_28),.acc(r1_28),.res(r1_29),.clk(clk),.wout(w1_29));
	PE pe1_30(.x(x30),.w(w1_29),.acc(r1_29),.res(r1_30),.clk(clk),.wout(w1_30));
	PE pe1_31(.x(x31),.w(w1_30),.acc(r1_30),.res(r1_31),.clk(clk),.wout(w1_31));
	PE pe1_32(.x(x32),.w(w1_31),.acc(r1_31),.res(r1_32),.clk(clk),.wout(w1_32));
	PE pe1_33(.x(x33),.w(w1_32),.acc(r1_32),.res(r1_33),.clk(clk),.wout(w1_33));
	PE pe1_34(.x(x34),.w(w1_33),.acc(r1_33),.res(r1_34),.clk(clk),.wout(w1_34));
	PE pe1_35(.x(x35),.w(w1_34),.acc(r1_34),.res(r1_35),.clk(clk),.wout(w1_35));
	PE pe1_36(.x(x36),.w(w1_35),.acc(r1_35),.res(r1_36),.clk(clk),.wout(w1_36));
	PE pe1_37(.x(x37),.w(w1_36),.acc(r1_36),.res(r1_37),.clk(clk),.wout(w1_37));
	PE pe1_38(.x(x38),.w(w1_37),.acc(r1_37),.res(r1_38),.clk(clk),.wout(w1_38));
	PE pe1_39(.x(x39),.w(w1_38),.acc(r1_38),.res(r1_39),.clk(clk),.wout(w1_39));
	PE pe1_40(.x(x40),.w(w1_39),.acc(r1_39),.res(r1_40),.clk(clk),.wout(w1_40));
	PE pe1_41(.x(x41),.w(w1_40),.acc(r1_40),.res(r1_41),.clk(clk),.wout(w1_41));
	PE pe1_42(.x(x42),.w(w1_41),.acc(r1_41),.res(r1_42),.clk(clk),.wout(w1_42));
	PE pe1_43(.x(x43),.w(w1_42),.acc(r1_42),.res(r1_43),.clk(clk),.wout(w1_43));
	PE pe1_44(.x(x44),.w(w1_43),.acc(r1_43),.res(r1_44),.clk(clk),.wout(w1_44));
	PE pe1_45(.x(x45),.w(w1_44),.acc(r1_44),.res(r1_45),.clk(clk),.wout(w1_45));
	PE pe1_46(.x(x46),.w(w1_45),.acc(r1_45),.res(r1_46),.clk(clk),.wout(w1_46));
	PE pe1_47(.x(x47),.w(w1_46),.acc(r1_46),.res(r1_47),.clk(clk),.wout(w1_47));
	PE pe1_48(.x(x48),.w(w1_47),.acc(r1_47),.res(r1_48),.clk(clk),.wout(w1_48));
	PE pe1_49(.x(x49),.w(w1_48),.acc(r1_48),.res(r1_49),.clk(clk),.wout(w1_49));
	PE pe1_50(.x(x50),.w(w1_49),.acc(r1_49),.res(r1_50),.clk(clk),.wout(w1_50));
	PE pe1_51(.x(x51),.w(w1_50),.acc(r1_50),.res(r1_51),.clk(clk),.wout(w1_51));
	PE pe1_52(.x(x52),.w(w1_51),.acc(r1_51),.res(r1_52),.clk(clk),.wout(w1_52));
	PE pe1_53(.x(x53),.w(w1_52),.acc(r1_52),.res(r1_53),.clk(clk),.wout(w1_53));
	PE pe1_54(.x(x54),.w(w1_53),.acc(r1_53),.res(r1_54),.clk(clk),.wout(w1_54));
	PE pe1_55(.x(x55),.w(w1_54),.acc(r1_54),.res(r1_55),.clk(clk),.wout(w1_55));
	PE pe1_56(.x(x56),.w(w1_55),.acc(r1_55),.res(r1_56),.clk(clk),.wout(w1_56));
	PE pe1_57(.x(x57),.w(w1_56),.acc(r1_56),.res(r1_57),.clk(clk),.wout(w1_57));
	PE pe1_58(.x(x58),.w(w1_57),.acc(r1_57),.res(r1_58),.clk(clk),.wout(w1_58));
	PE pe1_59(.x(x59),.w(w1_58),.acc(r1_58),.res(r1_59),.clk(clk),.wout(w1_59));
	PE pe1_60(.x(x60),.w(w1_59),.acc(r1_59),.res(r1_60),.clk(clk),.wout(w1_60));
	PE pe1_61(.x(x61),.w(w1_60),.acc(r1_60),.res(r1_61),.clk(clk),.wout(w1_61));
	PE pe1_62(.x(x62),.w(w1_61),.acc(r1_61),.res(r1_62),.clk(clk),.wout(w1_62));
	PE pe1_63(.x(x63),.w(w1_62),.acc(r1_62),.res(r1_63),.clk(clk),.wout(w1_63));
	PE pe1_64(.x(x64),.w(w1_63),.acc(r1_63),.res(r1_64),.clk(clk),.wout(w1_64));
	PE pe1_65(.x(x65),.w(w1_64),.acc(r1_64),.res(r1_65),.clk(clk),.wout(w1_65));
	PE pe1_66(.x(x66),.w(w1_65),.acc(r1_65),.res(r1_66),.clk(clk),.wout(w1_66));
	PE pe1_67(.x(x67),.w(w1_66),.acc(r1_66),.res(r1_67),.clk(clk),.wout(w1_67));
	PE pe1_68(.x(x68),.w(w1_67),.acc(r1_67),.res(r1_68),.clk(clk),.wout(w1_68));
	PE pe1_69(.x(x69),.w(w1_68),.acc(r1_68),.res(r1_69),.clk(clk),.wout(w1_69));
	PE pe1_70(.x(x70),.w(w1_69),.acc(r1_69),.res(r1_70),.clk(clk),.wout(w1_70));
	PE pe1_71(.x(x71),.w(w1_70),.acc(r1_70),.res(r1_71),.clk(clk),.wout(w1_71));
	PE pe1_72(.x(x72),.w(w1_71),.acc(r1_71),.res(r1_72),.clk(clk),.wout(w1_72));
	PE pe1_73(.x(x73),.w(w1_72),.acc(r1_72),.res(r1_73),.clk(clk),.wout(w1_73));
	PE pe1_74(.x(x74),.w(w1_73),.acc(r1_73),.res(r1_74),.clk(clk),.wout(w1_74));
	PE pe1_75(.x(x75),.w(w1_74),.acc(r1_74),.res(r1_75),.clk(clk),.wout(w1_75));
	PE pe1_76(.x(x76),.w(w1_75),.acc(r1_75),.res(r1_76),.clk(clk),.wout(w1_76));
	PE pe1_77(.x(x77),.w(w1_76),.acc(r1_76),.res(r1_77),.clk(clk),.wout(w1_77));
	PE pe1_78(.x(x78),.w(w1_77),.acc(r1_77),.res(r1_78),.clk(clk),.wout(w1_78));
	PE pe1_79(.x(x79),.w(w1_78),.acc(r1_78),.res(r1_79),.clk(clk),.wout(w1_79));
	PE pe1_80(.x(x80),.w(w1_79),.acc(r1_79),.res(r1_80),.clk(clk),.wout(w1_80));
	PE pe1_81(.x(x81),.w(w1_80),.acc(r1_80),.res(r1_81),.clk(clk),.wout(w1_81));
	PE pe1_82(.x(x82),.w(w1_81),.acc(r1_81),.res(r1_82),.clk(clk),.wout(w1_82));
	PE pe1_83(.x(x83),.w(w1_82),.acc(r1_82),.res(r1_83),.clk(clk),.wout(w1_83));
	PE pe1_84(.x(x84),.w(w1_83),.acc(r1_83),.res(r1_84),.clk(clk),.wout(w1_84));
	PE pe1_85(.x(x85),.w(w1_84),.acc(r1_84),.res(r1_85),.clk(clk),.wout(w1_85));
	PE pe1_86(.x(x86),.w(w1_85),.acc(r1_85),.res(r1_86),.clk(clk),.wout(w1_86));
	PE pe1_87(.x(x87),.w(w1_86),.acc(r1_86),.res(r1_87),.clk(clk),.wout(w1_87));
	PE pe1_88(.x(x88),.w(w1_87),.acc(r1_87),.res(r1_88),.clk(clk),.wout(w1_88));
	PE pe1_89(.x(x89),.w(w1_88),.acc(r1_88),.res(r1_89),.clk(clk),.wout(w1_89));
	PE pe1_90(.x(x90),.w(w1_89),.acc(r1_89),.res(r1_90),.clk(clk),.wout(w1_90));
	PE pe1_91(.x(x91),.w(w1_90),.acc(r1_90),.res(r1_91),.clk(clk),.wout(w1_91));
	PE pe1_92(.x(x92),.w(w1_91),.acc(r1_91),.res(r1_92),.clk(clk),.wout(w1_92));
	PE pe1_93(.x(x93),.w(w1_92),.acc(r1_92),.res(r1_93),.clk(clk),.wout(w1_93));
	PE pe1_94(.x(x94),.w(w1_93),.acc(r1_93),.res(r1_94),.clk(clk),.wout(w1_94));
	PE pe1_95(.x(x95),.w(w1_94),.acc(r1_94),.res(r1_95),.clk(clk),.wout(w1_95));
	PE pe1_96(.x(x96),.w(w1_95),.acc(r1_95),.res(r1_96),.clk(clk),.wout(w1_96));
	PE pe1_97(.x(x97),.w(w1_96),.acc(r1_96),.res(r1_97),.clk(clk),.wout(w1_97));
	PE pe1_98(.x(x98),.w(w1_97),.acc(r1_97),.res(r1_98),.clk(clk),.wout(w1_98));
	PE pe1_99(.x(x99),.w(w1_98),.acc(r1_98),.res(r1_99),.clk(clk),.wout(w1_99));
	PE pe1_100(.x(x100),.w(w1_99),.acc(r1_99),.res(r1_100),.clk(clk),.wout(w1_100));
	PE pe1_101(.x(x101),.w(w1_100),.acc(r1_100),.res(r1_101),.clk(clk),.wout(w1_101));
	PE pe1_102(.x(x102),.w(w1_101),.acc(r1_101),.res(r1_102),.clk(clk),.wout(w1_102));
	PE pe1_103(.x(x103),.w(w1_102),.acc(r1_102),.res(r1_103),.clk(clk),.wout(w1_103));
	PE pe1_104(.x(x104),.w(w1_103),.acc(r1_103),.res(r1_104),.clk(clk),.wout(w1_104));
	PE pe1_105(.x(x105),.w(w1_104),.acc(r1_104),.res(r1_105),.clk(clk),.wout(w1_105));
	PE pe1_106(.x(x106),.w(w1_105),.acc(r1_105),.res(r1_106),.clk(clk),.wout(w1_106));
	PE pe1_107(.x(x107),.w(w1_106),.acc(r1_106),.res(r1_107),.clk(clk),.wout(w1_107));
	PE pe1_108(.x(x108),.w(w1_107),.acc(r1_107),.res(r1_108),.clk(clk),.wout(w1_108));
	PE pe1_109(.x(x109),.w(w1_108),.acc(r1_108),.res(r1_109),.clk(clk),.wout(w1_109));
	PE pe1_110(.x(x110),.w(w1_109),.acc(r1_109),.res(r1_110),.clk(clk),.wout(w1_110));
	PE pe1_111(.x(x111),.w(w1_110),.acc(r1_110),.res(r1_111),.clk(clk),.wout(w1_111));
	PE pe1_112(.x(x112),.w(w1_111),.acc(r1_111),.res(r1_112),.clk(clk),.wout(w1_112));
	PE pe1_113(.x(x113),.w(w1_112),.acc(r1_112),.res(r1_113),.clk(clk),.wout(w1_113));
	PE pe1_114(.x(x114),.w(w1_113),.acc(r1_113),.res(r1_114),.clk(clk),.wout(w1_114));
	PE pe1_115(.x(x115),.w(w1_114),.acc(r1_114),.res(r1_115),.clk(clk),.wout(w1_115));
	PE pe1_116(.x(x116),.w(w1_115),.acc(r1_115),.res(r1_116),.clk(clk),.wout(w1_116));
	PE pe1_117(.x(x117),.w(w1_116),.acc(r1_116),.res(r1_117),.clk(clk),.wout(w1_117));
	PE pe1_118(.x(x118),.w(w1_117),.acc(r1_117),.res(r1_118),.clk(clk),.wout(w1_118));
	PE pe1_119(.x(x119),.w(w1_118),.acc(r1_118),.res(r1_119),.clk(clk),.wout(w1_119));
	PE pe1_120(.x(x120),.w(w1_119),.acc(r1_119),.res(r1_120),.clk(clk),.wout(w1_120));
	PE pe1_121(.x(x121),.w(w1_120),.acc(r1_120),.res(r1_121),.clk(clk),.wout(w1_121));
	PE pe1_122(.x(x122),.w(w1_121),.acc(r1_121),.res(r1_122),.clk(clk),.wout(w1_122));
	PE pe1_123(.x(x123),.w(w1_122),.acc(r1_122),.res(r1_123),.clk(clk),.wout(w1_123));
	PE pe1_124(.x(x124),.w(w1_123),.acc(r1_123),.res(r1_124),.clk(clk),.wout(w1_124));
	PE pe1_125(.x(x125),.w(w1_124),.acc(r1_124),.res(r1_125),.clk(clk),.wout(w1_125));
	PE pe1_126(.x(x126),.w(w1_125),.acc(r1_125),.res(r1_126),.clk(clk),.wout(w1_126));
	PE pe1_127(.x(x127),.w(w1_126),.acc(r1_126),.res(result1),.clk(clk),.wout(weight1));

	PE pe2_0(.x(x0),.w(w2),.acc(32'h0),.res(r2_0),.clk(clk),.wout(w2_0));
	PE pe2_1(.x(x1),.w(w2_0),.acc(r2_0),.res(r2_1),.clk(clk),.wout(w2_1));
	PE pe2_2(.x(x2),.w(w2_1),.acc(r2_1),.res(r2_2),.clk(clk),.wout(w2_2));
	PE pe2_3(.x(x3),.w(w2_2),.acc(r2_2),.res(r2_3),.clk(clk),.wout(w2_3));
	PE pe2_4(.x(x4),.w(w2_3),.acc(r2_3),.res(r2_4),.clk(clk),.wout(w2_4));
	PE pe2_5(.x(x5),.w(w2_4),.acc(r2_4),.res(r2_5),.clk(clk),.wout(w2_5));
	PE pe2_6(.x(x6),.w(w2_5),.acc(r2_5),.res(r2_6),.clk(clk),.wout(w2_6));
	PE pe2_7(.x(x7),.w(w2_6),.acc(r2_6),.res(r2_7),.clk(clk),.wout(w2_7));
	PE pe2_8(.x(x8),.w(w2_7),.acc(r2_7),.res(r2_8),.clk(clk),.wout(w2_8));
	PE pe2_9(.x(x9),.w(w2_8),.acc(r2_8),.res(r2_9),.clk(clk),.wout(w2_9));
	PE pe2_10(.x(x10),.w(w2_9),.acc(r2_9),.res(r2_10),.clk(clk),.wout(w2_10));
	PE pe2_11(.x(x11),.w(w2_10),.acc(r2_10),.res(r2_11),.clk(clk),.wout(w2_11));
	PE pe2_12(.x(x12),.w(w2_11),.acc(r2_11),.res(r2_12),.clk(clk),.wout(w2_12));
	PE pe2_13(.x(x13),.w(w2_12),.acc(r2_12),.res(r2_13),.clk(clk),.wout(w2_13));
	PE pe2_14(.x(x14),.w(w2_13),.acc(r2_13),.res(r2_14),.clk(clk),.wout(w2_14));
	PE pe2_15(.x(x15),.w(w2_14),.acc(r2_14),.res(r2_15),.clk(clk),.wout(w2_15));
	PE pe2_16(.x(x16),.w(w2_15),.acc(r2_15),.res(r2_16),.clk(clk),.wout(w2_16));
	PE pe2_17(.x(x17),.w(w2_16),.acc(r2_16),.res(r2_17),.clk(clk),.wout(w2_17));
	PE pe2_18(.x(x18),.w(w2_17),.acc(r2_17),.res(r2_18),.clk(clk),.wout(w2_18));
	PE pe2_19(.x(x19),.w(w2_18),.acc(r2_18),.res(r2_19),.clk(clk),.wout(w2_19));
	PE pe2_20(.x(x20),.w(w2_19),.acc(r2_19),.res(r2_20),.clk(clk),.wout(w2_20));
	PE pe2_21(.x(x21),.w(w2_20),.acc(r2_20),.res(r2_21),.clk(clk),.wout(w2_21));
	PE pe2_22(.x(x22),.w(w2_21),.acc(r2_21),.res(r2_22),.clk(clk),.wout(w2_22));
	PE pe2_23(.x(x23),.w(w2_22),.acc(r2_22),.res(r2_23),.clk(clk),.wout(w2_23));
	PE pe2_24(.x(x24),.w(w2_23),.acc(r2_23),.res(r2_24),.clk(clk),.wout(w2_24));
	PE pe2_25(.x(x25),.w(w2_24),.acc(r2_24),.res(r2_25),.clk(clk),.wout(w2_25));
	PE pe2_26(.x(x26),.w(w2_25),.acc(r2_25),.res(r2_26),.clk(clk),.wout(w2_26));
	PE pe2_27(.x(x27),.w(w2_26),.acc(r2_26),.res(r2_27),.clk(clk),.wout(w2_27));
	PE pe2_28(.x(x28),.w(w2_27),.acc(r2_27),.res(r2_28),.clk(clk),.wout(w2_28));
	PE pe2_29(.x(x29),.w(w2_28),.acc(r2_28),.res(r2_29),.clk(clk),.wout(w2_29));
	PE pe2_30(.x(x30),.w(w2_29),.acc(r2_29),.res(r2_30),.clk(clk),.wout(w2_30));
	PE pe2_31(.x(x31),.w(w2_30),.acc(r2_30),.res(r2_31),.clk(clk),.wout(w2_31));
	PE pe2_32(.x(x32),.w(w2_31),.acc(r2_31),.res(r2_32),.clk(clk),.wout(w2_32));
	PE pe2_33(.x(x33),.w(w2_32),.acc(r2_32),.res(r2_33),.clk(clk),.wout(w2_33));
	PE pe2_34(.x(x34),.w(w2_33),.acc(r2_33),.res(r2_34),.clk(clk),.wout(w2_34));
	PE pe2_35(.x(x35),.w(w2_34),.acc(r2_34),.res(r2_35),.clk(clk),.wout(w2_35));
	PE pe2_36(.x(x36),.w(w2_35),.acc(r2_35),.res(r2_36),.clk(clk),.wout(w2_36));
	PE pe2_37(.x(x37),.w(w2_36),.acc(r2_36),.res(r2_37),.clk(clk),.wout(w2_37));
	PE pe2_38(.x(x38),.w(w2_37),.acc(r2_37),.res(r2_38),.clk(clk),.wout(w2_38));
	PE pe2_39(.x(x39),.w(w2_38),.acc(r2_38),.res(r2_39),.clk(clk),.wout(w2_39));
	PE pe2_40(.x(x40),.w(w2_39),.acc(r2_39),.res(r2_40),.clk(clk),.wout(w2_40));
	PE pe2_41(.x(x41),.w(w2_40),.acc(r2_40),.res(r2_41),.clk(clk),.wout(w2_41));
	PE pe2_42(.x(x42),.w(w2_41),.acc(r2_41),.res(r2_42),.clk(clk),.wout(w2_42));
	PE pe2_43(.x(x43),.w(w2_42),.acc(r2_42),.res(r2_43),.clk(clk),.wout(w2_43));
	PE pe2_44(.x(x44),.w(w2_43),.acc(r2_43),.res(r2_44),.clk(clk),.wout(w2_44));
	PE pe2_45(.x(x45),.w(w2_44),.acc(r2_44),.res(r2_45),.clk(clk),.wout(w2_45));
	PE pe2_46(.x(x46),.w(w2_45),.acc(r2_45),.res(r2_46),.clk(clk),.wout(w2_46));
	PE pe2_47(.x(x47),.w(w2_46),.acc(r2_46),.res(r2_47),.clk(clk),.wout(w2_47));
	PE pe2_48(.x(x48),.w(w2_47),.acc(r2_47),.res(r2_48),.clk(clk),.wout(w2_48));
	PE pe2_49(.x(x49),.w(w2_48),.acc(r2_48),.res(r2_49),.clk(clk),.wout(w2_49));
	PE pe2_50(.x(x50),.w(w2_49),.acc(r2_49),.res(r2_50),.clk(clk),.wout(w2_50));
	PE pe2_51(.x(x51),.w(w2_50),.acc(r2_50),.res(r2_51),.clk(clk),.wout(w2_51));
	PE pe2_52(.x(x52),.w(w2_51),.acc(r2_51),.res(r2_52),.clk(clk),.wout(w2_52));
	PE pe2_53(.x(x53),.w(w2_52),.acc(r2_52),.res(r2_53),.clk(clk),.wout(w2_53));
	PE pe2_54(.x(x54),.w(w2_53),.acc(r2_53),.res(r2_54),.clk(clk),.wout(w2_54));
	PE pe2_55(.x(x55),.w(w2_54),.acc(r2_54),.res(r2_55),.clk(clk),.wout(w2_55));
	PE pe2_56(.x(x56),.w(w2_55),.acc(r2_55),.res(r2_56),.clk(clk),.wout(w2_56));
	PE pe2_57(.x(x57),.w(w2_56),.acc(r2_56),.res(r2_57),.clk(clk),.wout(w2_57));
	PE pe2_58(.x(x58),.w(w2_57),.acc(r2_57),.res(r2_58),.clk(clk),.wout(w2_58));
	PE pe2_59(.x(x59),.w(w2_58),.acc(r2_58),.res(r2_59),.clk(clk),.wout(w2_59));
	PE pe2_60(.x(x60),.w(w2_59),.acc(r2_59),.res(r2_60),.clk(clk),.wout(w2_60));
	PE pe2_61(.x(x61),.w(w2_60),.acc(r2_60),.res(r2_61),.clk(clk),.wout(w2_61));
	PE pe2_62(.x(x62),.w(w2_61),.acc(r2_61),.res(r2_62),.clk(clk),.wout(w2_62));
	PE pe2_63(.x(x63),.w(w2_62),.acc(r2_62),.res(r2_63),.clk(clk),.wout(w2_63));
	PE pe2_64(.x(x64),.w(w2_63),.acc(r2_63),.res(r2_64),.clk(clk),.wout(w2_64));
	PE pe2_65(.x(x65),.w(w2_64),.acc(r2_64),.res(r2_65),.clk(clk),.wout(w2_65));
	PE pe2_66(.x(x66),.w(w2_65),.acc(r2_65),.res(r2_66),.clk(clk),.wout(w2_66));
	PE pe2_67(.x(x67),.w(w2_66),.acc(r2_66),.res(r2_67),.clk(clk),.wout(w2_67));
	PE pe2_68(.x(x68),.w(w2_67),.acc(r2_67),.res(r2_68),.clk(clk),.wout(w2_68));
	PE pe2_69(.x(x69),.w(w2_68),.acc(r2_68),.res(r2_69),.clk(clk),.wout(w2_69));
	PE pe2_70(.x(x70),.w(w2_69),.acc(r2_69),.res(r2_70),.clk(clk),.wout(w2_70));
	PE pe2_71(.x(x71),.w(w2_70),.acc(r2_70),.res(r2_71),.clk(clk),.wout(w2_71));
	PE pe2_72(.x(x72),.w(w2_71),.acc(r2_71),.res(r2_72),.clk(clk),.wout(w2_72));
	PE pe2_73(.x(x73),.w(w2_72),.acc(r2_72),.res(r2_73),.clk(clk),.wout(w2_73));
	PE pe2_74(.x(x74),.w(w2_73),.acc(r2_73),.res(r2_74),.clk(clk),.wout(w2_74));
	PE pe2_75(.x(x75),.w(w2_74),.acc(r2_74),.res(r2_75),.clk(clk),.wout(w2_75));
	PE pe2_76(.x(x76),.w(w2_75),.acc(r2_75),.res(r2_76),.clk(clk),.wout(w2_76));
	PE pe2_77(.x(x77),.w(w2_76),.acc(r2_76),.res(r2_77),.clk(clk),.wout(w2_77));
	PE pe2_78(.x(x78),.w(w2_77),.acc(r2_77),.res(r2_78),.clk(clk),.wout(w2_78));
	PE pe2_79(.x(x79),.w(w2_78),.acc(r2_78),.res(r2_79),.clk(clk),.wout(w2_79));
	PE pe2_80(.x(x80),.w(w2_79),.acc(r2_79),.res(r2_80),.clk(clk),.wout(w2_80));
	PE pe2_81(.x(x81),.w(w2_80),.acc(r2_80),.res(r2_81),.clk(clk),.wout(w2_81));
	PE pe2_82(.x(x82),.w(w2_81),.acc(r2_81),.res(r2_82),.clk(clk),.wout(w2_82));
	PE pe2_83(.x(x83),.w(w2_82),.acc(r2_82),.res(r2_83),.clk(clk),.wout(w2_83));
	PE pe2_84(.x(x84),.w(w2_83),.acc(r2_83),.res(r2_84),.clk(clk),.wout(w2_84));
	PE pe2_85(.x(x85),.w(w2_84),.acc(r2_84),.res(r2_85),.clk(clk),.wout(w2_85));
	PE pe2_86(.x(x86),.w(w2_85),.acc(r2_85),.res(r2_86),.clk(clk),.wout(w2_86));
	PE pe2_87(.x(x87),.w(w2_86),.acc(r2_86),.res(r2_87),.clk(clk),.wout(w2_87));
	PE pe2_88(.x(x88),.w(w2_87),.acc(r2_87),.res(r2_88),.clk(clk),.wout(w2_88));
	PE pe2_89(.x(x89),.w(w2_88),.acc(r2_88),.res(r2_89),.clk(clk),.wout(w2_89));
	PE pe2_90(.x(x90),.w(w2_89),.acc(r2_89),.res(r2_90),.clk(clk),.wout(w2_90));
	PE pe2_91(.x(x91),.w(w2_90),.acc(r2_90),.res(r2_91),.clk(clk),.wout(w2_91));
	PE pe2_92(.x(x92),.w(w2_91),.acc(r2_91),.res(r2_92),.clk(clk),.wout(w2_92));
	PE pe2_93(.x(x93),.w(w2_92),.acc(r2_92),.res(r2_93),.clk(clk),.wout(w2_93));
	PE pe2_94(.x(x94),.w(w2_93),.acc(r2_93),.res(r2_94),.clk(clk),.wout(w2_94));
	PE pe2_95(.x(x95),.w(w2_94),.acc(r2_94),.res(r2_95),.clk(clk),.wout(w2_95));
	PE pe2_96(.x(x96),.w(w2_95),.acc(r2_95),.res(r2_96),.clk(clk),.wout(w2_96));
	PE pe2_97(.x(x97),.w(w2_96),.acc(r2_96),.res(r2_97),.clk(clk),.wout(w2_97));
	PE pe2_98(.x(x98),.w(w2_97),.acc(r2_97),.res(r2_98),.clk(clk),.wout(w2_98));
	PE pe2_99(.x(x99),.w(w2_98),.acc(r2_98),.res(r2_99),.clk(clk),.wout(w2_99));
	PE pe2_100(.x(x100),.w(w2_99),.acc(r2_99),.res(r2_100),.clk(clk),.wout(w2_100));
	PE pe2_101(.x(x101),.w(w2_100),.acc(r2_100),.res(r2_101),.clk(clk),.wout(w2_101));
	PE pe2_102(.x(x102),.w(w2_101),.acc(r2_101),.res(r2_102),.clk(clk),.wout(w2_102));
	PE pe2_103(.x(x103),.w(w2_102),.acc(r2_102),.res(r2_103),.clk(clk),.wout(w2_103));
	PE pe2_104(.x(x104),.w(w2_103),.acc(r2_103),.res(r2_104),.clk(clk),.wout(w2_104));
	PE pe2_105(.x(x105),.w(w2_104),.acc(r2_104),.res(r2_105),.clk(clk),.wout(w2_105));
	PE pe2_106(.x(x106),.w(w2_105),.acc(r2_105),.res(r2_106),.clk(clk),.wout(w2_106));
	PE pe2_107(.x(x107),.w(w2_106),.acc(r2_106),.res(r2_107),.clk(clk),.wout(w2_107));
	PE pe2_108(.x(x108),.w(w2_107),.acc(r2_107),.res(r2_108),.clk(clk),.wout(w2_108));
	PE pe2_109(.x(x109),.w(w2_108),.acc(r2_108),.res(r2_109),.clk(clk),.wout(w2_109));
	PE pe2_110(.x(x110),.w(w2_109),.acc(r2_109),.res(r2_110),.clk(clk),.wout(w2_110));
	PE pe2_111(.x(x111),.w(w2_110),.acc(r2_110),.res(r2_111),.clk(clk),.wout(w2_111));
	PE pe2_112(.x(x112),.w(w2_111),.acc(r2_111),.res(r2_112),.clk(clk),.wout(w2_112));
	PE pe2_113(.x(x113),.w(w2_112),.acc(r2_112),.res(r2_113),.clk(clk),.wout(w2_113));
	PE pe2_114(.x(x114),.w(w2_113),.acc(r2_113),.res(r2_114),.clk(clk),.wout(w2_114));
	PE pe2_115(.x(x115),.w(w2_114),.acc(r2_114),.res(r2_115),.clk(clk),.wout(w2_115));
	PE pe2_116(.x(x116),.w(w2_115),.acc(r2_115),.res(r2_116),.clk(clk),.wout(w2_116));
	PE pe2_117(.x(x117),.w(w2_116),.acc(r2_116),.res(r2_117),.clk(clk),.wout(w2_117));
	PE pe2_118(.x(x118),.w(w2_117),.acc(r2_117),.res(r2_118),.clk(clk),.wout(w2_118));
	PE pe2_119(.x(x119),.w(w2_118),.acc(r2_118),.res(r2_119),.clk(clk),.wout(w2_119));
	PE pe2_120(.x(x120),.w(w2_119),.acc(r2_119),.res(r2_120),.clk(clk),.wout(w2_120));
	PE pe2_121(.x(x121),.w(w2_120),.acc(r2_120),.res(r2_121),.clk(clk),.wout(w2_121));
	PE pe2_122(.x(x122),.w(w2_121),.acc(r2_121),.res(r2_122),.clk(clk),.wout(w2_122));
	PE pe2_123(.x(x123),.w(w2_122),.acc(r2_122),.res(r2_123),.clk(clk),.wout(w2_123));
	PE pe2_124(.x(x124),.w(w2_123),.acc(r2_123),.res(r2_124),.clk(clk),.wout(w2_124));
	PE pe2_125(.x(x125),.w(w2_124),.acc(r2_124),.res(r2_125),.clk(clk),.wout(w2_125));
	PE pe2_126(.x(x126),.w(w2_125),.acc(r2_125),.res(r2_126),.clk(clk),.wout(w2_126));
	PE pe2_127(.x(x127),.w(w2_126),.acc(r2_126),.res(result2),.clk(clk),.wout(weight2));

	PE pe3_0(.x(x0),.w(w3),.acc(32'h0),.res(r3_0),.clk(clk),.wout(w3_0));
	PE pe3_1(.x(x1),.w(w3_0),.acc(r3_0),.res(r3_1),.clk(clk),.wout(w3_1));
	PE pe3_2(.x(x2),.w(w3_1),.acc(r3_1),.res(r3_2),.clk(clk),.wout(w3_2));
	PE pe3_3(.x(x3),.w(w3_2),.acc(r3_2),.res(r3_3),.clk(clk),.wout(w3_3));
	PE pe3_4(.x(x4),.w(w3_3),.acc(r3_3),.res(r3_4),.clk(clk),.wout(w3_4));
	PE pe3_5(.x(x5),.w(w3_4),.acc(r3_4),.res(r3_5),.clk(clk),.wout(w3_5));
	PE pe3_6(.x(x6),.w(w3_5),.acc(r3_5),.res(r3_6),.clk(clk),.wout(w3_6));
	PE pe3_7(.x(x7),.w(w3_6),.acc(r3_6),.res(r3_7),.clk(clk),.wout(w3_7));
	PE pe3_8(.x(x8),.w(w3_7),.acc(r3_7),.res(r3_8),.clk(clk),.wout(w3_8));
	PE pe3_9(.x(x9),.w(w3_8),.acc(r3_8),.res(r3_9),.clk(clk),.wout(w3_9));
	PE pe3_10(.x(x10),.w(w3_9),.acc(r3_9),.res(r3_10),.clk(clk),.wout(w3_10));
	PE pe3_11(.x(x11),.w(w3_10),.acc(r3_10),.res(r3_11),.clk(clk),.wout(w3_11));
	PE pe3_12(.x(x12),.w(w3_11),.acc(r3_11),.res(r3_12),.clk(clk),.wout(w3_12));
	PE pe3_13(.x(x13),.w(w3_12),.acc(r3_12),.res(r3_13),.clk(clk),.wout(w3_13));
	PE pe3_14(.x(x14),.w(w3_13),.acc(r3_13),.res(r3_14),.clk(clk),.wout(w3_14));
	PE pe3_15(.x(x15),.w(w3_14),.acc(r3_14),.res(r3_15),.clk(clk),.wout(w3_15));
	PE pe3_16(.x(x16),.w(w3_15),.acc(r3_15),.res(r3_16),.clk(clk),.wout(w3_16));
	PE pe3_17(.x(x17),.w(w3_16),.acc(r3_16),.res(r3_17),.clk(clk),.wout(w3_17));
	PE pe3_18(.x(x18),.w(w3_17),.acc(r3_17),.res(r3_18),.clk(clk),.wout(w3_18));
	PE pe3_19(.x(x19),.w(w3_18),.acc(r3_18),.res(r3_19),.clk(clk),.wout(w3_19));
	PE pe3_20(.x(x20),.w(w3_19),.acc(r3_19),.res(r3_20),.clk(clk),.wout(w3_20));
	PE pe3_21(.x(x21),.w(w3_20),.acc(r3_20),.res(r3_21),.clk(clk),.wout(w3_21));
	PE pe3_22(.x(x22),.w(w3_21),.acc(r3_21),.res(r3_22),.clk(clk),.wout(w3_22));
	PE pe3_23(.x(x23),.w(w3_22),.acc(r3_22),.res(r3_23),.clk(clk),.wout(w3_23));
	PE pe3_24(.x(x24),.w(w3_23),.acc(r3_23),.res(r3_24),.clk(clk),.wout(w3_24));
	PE pe3_25(.x(x25),.w(w3_24),.acc(r3_24),.res(r3_25),.clk(clk),.wout(w3_25));
	PE pe3_26(.x(x26),.w(w3_25),.acc(r3_25),.res(r3_26),.clk(clk),.wout(w3_26));
	PE pe3_27(.x(x27),.w(w3_26),.acc(r3_26),.res(r3_27),.clk(clk),.wout(w3_27));
	PE pe3_28(.x(x28),.w(w3_27),.acc(r3_27),.res(r3_28),.clk(clk),.wout(w3_28));
	PE pe3_29(.x(x29),.w(w3_28),.acc(r3_28),.res(r3_29),.clk(clk),.wout(w3_29));
	PE pe3_30(.x(x30),.w(w3_29),.acc(r3_29),.res(r3_30),.clk(clk),.wout(w3_30));
	PE pe3_31(.x(x31),.w(w3_30),.acc(r3_30),.res(r3_31),.clk(clk),.wout(w3_31));
	PE pe3_32(.x(x32),.w(w3_31),.acc(r3_31),.res(r3_32),.clk(clk),.wout(w3_32));
	PE pe3_33(.x(x33),.w(w3_32),.acc(r3_32),.res(r3_33),.clk(clk),.wout(w3_33));
	PE pe3_34(.x(x34),.w(w3_33),.acc(r3_33),.res(r3_34),.clk(clk),.wout(w3_34));
	PE pe3_35(.x(x35),.w(w3_34),.acc(r3_34),.res(r3_35),.clk(clk),.wout(w3_35));
	PE pe3_36(.x(x36),.w(w3_35),.acc(r3_35),.res(r3_36),.clk(clk),.wout(w3_36));
	PE pe3_37(.x(x37),.w(w3_36),.acc(r3_36),.res(r3_37),.clk(clk),.wout(w3_37));
	PE pe3_38(.x(x38),.w(w3_37),.acc(r3_37),.res(r3_38),.clk(clk),.wout(w3_38));
	PE pe3_39(.x(x39),.w(w3_38),.acc(r3_38),.res(r3_39),.clk(clk),.wout(w3_39));
	PE pe3_40(.x(x40),.w(w3_39),.acc(r3_39),.res(r3_40),.clk(clk),.wout(w3_40));
	PE pe3_41(.x(x41),.w(w3_40),.acc(r3_40),.res(r3_41),.clk(clk),.wout(w3_41));
	PE pe3_42(.x(x42),.w(w3_41),.acc(r3_41),.res(r3_42),.clk(clk),.wout(w3_42));
	PE pe3_43(.x(x43),.w(w3_42),.acc(r3_42),.res(r3_43),.clk(clk),.wout(w3_43));
	PE pe3_44(.x(x44),.w(w3_43),.acc(r3_43),.res(r3_44),.clk(clk),.wout(w3_44));
	PE pe3_45(.x(x45),.w(w3_44),.acc(r3_44),.res(r3_45),.clk(clk),.wout(w3_45));
	PE pe3_46(.x(x46),.w(w3_45),.acc(r3_45),.res(r3_46),.clk(clk),.wout(w3_46));
	PE pe3_47(.x(x47),.w(w3_46),.acc(r3_46),.res(r3_47),.clk(clk),.wout(w3_47));
	PE pe3_48(.x(x48),.w(w3_47),.acc(r3_47),.res(r3_48),.clk(clk),.wout(w3_48));
	PE pe3_49(.x(x49),.w(w3_48),.acc(r3_48),.res(r3_49),.clk(clk),.wout(w3_49));
	PE pe3_50(.x(x50),.w(w3_49),.acc(r3_49),.res(r3_50),.clk(clk),.wout(w3_50));
	PE pe3_51(.x(x51),.w(w3_50),.acc(r3_50),.res(r3_51),.clk(clk),.wout(w3_51));
	PE pe3_52(.x(x52),.w(w3_51),.acc(r3_51),.res(r3_52),.clk(clk),.wout(w3_52));
	PE pe3_53(.x(x53),.w(w3_52),.acc(r3_52),.res(r3_53),.clk(clk),.wout(w3_53));
	PE pe3_54(.x(x54),.w(w3_53),.acc(r3_53),.res(r3_54),.clk(clk),.wout(w3_54));
	PE pe3_55(.x(x55),.w(w3_54),.acc(r3_54),.res(r3_55),.clk(clk),.wout(w3_55));
	PE pe3_56(.x(x56),.w(w3_55),.acc(r3_55),.res(r3_56),.clk(clk),.wout(w3_56));
	PE pe3_57(.x(x57),.w(w3_56),.acc(r3_56),.res(r3_57),.clk(clk),.wout(w3_57));
	PE pe3_58(.x(x58),.w(w3_57),.acc(r3_57),.res(r3_58),.clk(clk),.wout(w3_58));
	PE pe3_59(.x(x59),.w(w3_58),.acc(r3_58),.res(r3_59),.clk(clk),.wout(w3_59));
	PE pe3_60(.x(x60),.w(w3_59),.acc(r3_59),.res(r3_60),.clk(clk),.wout(w3_60));
	PE pe3_61(.x(x61),.w(w3_60),.acc(r3_60),.res(r3_61),.clk(clk),.wout(w3_61));
	PE pe3_62(.x(x62),.w(w3_61),.acc(r3_61),.res(r3_62),.clk(clk),.wout(w3_62));
	PE pe3_63(.x(x63),.w(w3_62),.acc(r3_62),.res(r3_63),.clk(clk),.wout(w3_63));
	PE pe3_64(.x(x64),.w(w3_63),.acc(r3_63),.res(r3_64),.clk(clk),.wout(w3_64));
	PE pe3_65(.x(x65),.w(w3_64),.acc(r3_64),.res(r3_65),.clk(clk),.wout(w3_65));
	PE pe3_66(.x(x66),.w(w3_65),.acc(r3_65),.res(r3_66),.clk(clk),.wout(w3_66));
	PE pe3_67(.x(x67),.w(w3_66),.acc(r3_66),.res(r3_67),.clk(clk),.wout(w3_67));
	PE pe3_68(.x(x68),.w(w3_67),.acc(r3_67),.res(r3_68),.clk(clk),.wout(w3_68));
	PE pe3_69(.x(x69),.w(w3_68),.acc(r3_68),.res(r3_69),.clk(clk),.wout(w3_69));
	PE pe3_70(.x(x70),.w(w3_69),.acc(r3_69),.res(r3_70),.clk(clk),.wout(w3_70));
	PE pe3_71(.x(x71),.w(w3_70),.acc(r3_70),.res(r3_71),.clk(clk),.wout(w3_71));
	PE pe3_72(.x(x72),.w(w3_71),.acc(r3_71),.res(r3_72),.clk(clk),.wout(w3_72));
	PE pe3_73(.x(x73),.w(w3_72),.acc(r3_72),.res(r3_73),.clk(clk),.wout(w3_73));
	PE pe3_74(.x(x74),.w(w3_73),.acc(r3_73),.res(r3_74),.clk(clk),.wout(w3_74));
	PE pe3_75(.x(x75),.w(w3_74),.acc(r3_74),.res(r3_75),.clk(clk),.wout(w3_75));
	PE pe3_76(.x(x76),.w(w3_75),.acc(r3_75),.res(r3_76),.clk(clk),.wout(w3_76));
	PE pe3_77(.x(x77),.w(w3_76),.acc(r3_76),.res(r3_77),.clk(clk),.wout(w3_77));
	PE pe3_78(.x(x78),.w(w3_77),.acc(r3_77),.res(r3_78),.clk(clk),.wout(w3_78));
	PE pe3_79(.x(x79),.w(w3_78),.acc(r3_78),.res(r3_79),.clk(clk),.wout(w3_79));
	PE pe3_80(.x(x80),.w(w3_79),.acc(r3_79),.res(r3_80),.clk(clk),.wout(w3_80));
	PE pe3_81(.x(x81),.w(w3_80),.acc(r3_80),.res(r3_81),.clk(clk),.wout(w3_81));
	PE pe3_82(.x(x82),.w(w3_81),.acc(r3_81),.res(r3_82),.clk(clk),.wout(w3_82));
	PE pe3_83(.x(x83),.w(w3_82),.acc(r3_82),.res(r3_83),.clk(clk),.wout(w3_83));
	PE pe3_84(.x(x84),.w(w3_83),.acc(r3_83),.res(r3_84),.clk(clk),.wout(w3_84));
	PE pe3_85(.x(x85),.w(w3_84),.acc(r3_84),.res(r3_85),.clk(clk),.wout(w3_85));
	PE pe3_86(.x(x86),.w(w3_85),.acc(r3_85),.res(r3_86),.clk(clk),.wout(w3_86));
	PE pe3_87(.x(x87),.w(w3_86),.acc(r3_86),.res(r3_87),.clk(clk),.wout(w3_87));
	PE pe3_88(.x(x88),.w(w3_87),.acc(r3_87),.res(r3_88),.clk(clk),.wout(w3_88));
	PE pe3_89(.x(x89),.w(w3_88),.acc(r3_88),.res(r3_89),.clk(clk),.wout(w3_89));
	PE pe3_90(.x(x90),.w(w3_89),.acc(r3_89),.res(r3_90),.clk(clk),.wout(w3_90));
	PE pe3_91(.x(x91),.w(w3_90),.acc(r3_90),.res(r3_91),.clk(clk),.wout(w3_91));
	PE pe3_92(.x(x92),.w(w3_91),.acc(r3_91),.res(r3_92),.clk(clk),.wout(w3_92));
	PE pe3_93(.x(x93),.w(w3_92),.acc(r3_92),.res(r3_93),.clk(clk),.wout(w3_93));
	PE pe3_94(.x(x94),.w(w3_93),.acc(r3_93),.res(r3_94),.clk(clk),.wout(w3_94));
	PE pe3_95(.x(x95),.w(w3_94),.acc(r3_94),.res(r3_95),.clk(clk),.wout(w3_95));
	PE pe3_96(.x(x96),.w(w3_95),.acc(r3_95),.res(r3_96),.clk(clk),.wout(w3_96));
	PE pe3_97(.x(x97),.w(w3_96),.acc(r3_96),.res(r3_97),.clk(clk),.wout(w3_97));
	PE pe3_98(.x(x98),.w(w3_97),.acc(r3_97),.res(r3_98),.clk(clk),.wout(w3_98));
	PE pe3_99(.x(x99),.w(w3_98),.acc(r3_98),.res(r3_99),.clk(clk),.wout(w3_99));
	PE pe3_100(.x(x100),.w(w3_99),.acc(r3_99),.res(r3_100),.clk(clk),.wout(w3_100));
	PE pe3_101(.x(x101),.w(w3_100),.acc(r3_100),.res(r3_101),.clk(clk),.wout(w3_101));
	PE pe3_102(.x(x102),.w(w3_101),.acc(r3_101),.res(r3_102),.clk(clk),.wout(w3_102));
	PE pe3_103(.x(x103),.w(w3_102),.acc(r3_102),.res(r3_103),.clk(clk),.wout(w3_103));
	PE pe3_104(.x(x104),.w(w3_103),.acc(r3_103),.res(r3_104),.clk(clk),.wout(w3_104));
	PE pe3_105(.x(x105),.w(w3_104),.acc(r3_104),.res(r3_105),.clk(clk),.wout(w3_105));
	PE pe3_106(.x(x106),.w(w3_105),.acc(r3_105),.res(r3_106),.clk(clk),.wout(w3_106));
	PE pe3_107(.x(x107),.w(w3_106),.acc(r3_106),.res(r3_107),.clk(clk),.wout(w3_107));
	PE pe3_108(.x(x108),.w(w3_107),.acc(r3_107),.res(r3_108),.clk(clk),.wout(w3_108));
	PE pe3_109(.x(x109),.w(w3_108),.acc(r3_108),.res(r3_109),.clk(clk),.wout(w3_109));
	PE pe3_110(.x(x110),.w(w3_109),.acc(r3_109),.res(r3_110),.clk(clk),.wout(w3_110));
	PE pe3_111(.x(x111),.w(w3_110),.acc(r3_110),.res(r3_111),.clk(clk),.wout(w3_111));
	PE pe3_112(.x(x112),.w(w3_111),.acc(r3_111),.res(r3_112),.clk(clk),.wout(w3_112));
	PE pe3_113(.x(x113),.w(w3_112),.acc(r3_112),.res(r3_113),.clk(clk),.wout(w3_113));
	PE pe3_114(.x(x114),.w(w3_113),.acc(r3_113),.res(r3_114),.clk(clk),.wout(w3_114));
	PE pe3_115(.x(x115),.w(w3_114),.acc(r3_114),.res(r3_115),.clk(clk),.wout(w3_115));
	PE pe3_116(.x(x116),.w(w3_115),.acc(r3_115),.res(r3_116),.clk(clk),.wout(w3_116));
	PE pe3_117(.x(x117),.w(w3_116),.acc(r3_116),.res(r3_117),.clk(clk),.wout(w3_117));
	PE pe3_118(.x(x118),.w(w3_117),.acc(r3_117),.res(r3_118),.clk(clk),.wout(w3_118));
	PE pe3_119(.x(x119),.w(w3_118),.acc(r3_118),.res(r3_119),.clk(clk),.wout(w3_119));
	PE pe3_120(.x(x120),.w(w3_119),.acc(r3_119),.res(r3_120),.clk(clk),.wout(w3_120));
	PE pe3_121(.x(x121),.w(w3_120),.acc(r3_120),.res(r3_121),.clk(clk),.wout(w3_121));
	PE pe3_122(.x(x122),.w(w3_121),.acc(r3_121),.res(r3_122),.clk(clk),.wout(w3_122));
	PE pe3_123(.x(x123),.w(w3_122),.acc(r3_122),.res(r3_123),.clk(clk),.wout(w3_123));
	PE pe3_124(.x(x124),.w(w3_123),.acc(r3_123),.res(r3_124),.clk(clk),.wout(w3_124));
	PE pe3_125(.x(x125),.w(w3_124),.acc(r3_124),.res(r3_125),.clk(clk),.wout(w3_125));
	PE pe3_126(.x(x126),.w(w3_125),.acc(r3_125),.res(r3_126),.clk(clk),.wout(w3_126));
	PE pe3_127(.x(x127),.w(w3_126),.acc(r3_126),.res(result3),.clk(clk),.wout(weight3));

	PE pe4_0(.x(x0),.w(w4),.acc(32'h0),.res(r4_0),.clk(clk),.wout(w4_0));
	PE pe4_1(.x(x1),.w(w4_0),.acc(r4_0),.res(r4_1),.clk(clk),.wout(w4_1));
	PE pe4_2(.x(x2),.w(w4_1),.acc(r4_1),.res(r4_2),.clk(clk),.wout(w4_2));
	PE pe4_3(.x(x3),.w(w4_2),.acc(r4_2),.res(r4_3),.clk(clk),.wout(w4_3));
	PE pe4_4(.x(x4),.w(w4_3),.acc(r4_3),.res(r4_4),.clk(clk),.wout(w4_4));
	PE pe4_5(.x(x5),.w(w4_4),.acc(r4_4),.res(r4_5),.clk(clk),.wout(w4_5));
	PE pe4_6(.x(x6),.w(w4_5),.acc(r4_5),.res(r4_6),.clk(clk),.wout(w4_6));
	PE pe4_7(.x(x7),.w(w4_6),.acc(r4_6),.res(r4_7),.clk(clk),.wout(w4_7));
	PE pe4_8(.x(x8),.w(w4_7),.acc(r4_7),.res(r4_8),.clk(clk),.wout(w4_8));
	PE pe4_9(.x(x9),.w(w4_8),.acc(r4_8),.res(r4_9),.clk(clk),.wout(w4_9));
	PE pe4_10(.x(x10),.w(w4_9),.acc(r4_9),.res(r4_10),.clk(clk),.wout(w4_10));
	PE pe4_11(.x(x11),.w(w4_10),.acc(r4_10),.res(r4_11),.clk(clk),.wout(w4_11));
	PE pe4_12(.x(x12),.w(w4_11),.acc(r4_11),.res(r4_12),.clk(clk),.wout(w4_12));
	PE pe4_13(.x(x13),.w(w4_12),.acc(r4_12),.res(r4_13),.clk(clk),.wout(w4_13));
	PE pe4_14(.x(x14),.w(w4_13),.acc(r4_13),.res(r4_14),.clk(clk),.wout(w4_14));
	PE pe4_15(.x(x15),.w(w4_14),.acc(r4_14),.res(r4_15),.clk(clk),.wout(w4_15));
	PE pe4_16(.x(x16),.w(w4_15),.acc(r4_15),.res(r4_16),.clk(clk),.wout(w4_16));
	PE pe4_17(.x(x17),.w(w4_16),.acc(r4_16),.res(r4_17),.clk(clk),.wout(w4_17));
	PE pe4_18(.x(x18),.w(w4_17),.acc(r4_17),.res(r4_18),.clk(clk),.wout(w4_18));
	PE pe4_19(.x(x19),.w(w4_18),.acc(r4_18),.res(r4_19),.clk(clk),.wout(w4_19));
	PE pe4_20(.x(x20),.w(w4_19),.acc(r4_19),.res(r4_20),.clk(clk),.wout(w4_20));
	PE pe4_21(.x(x21),.w(w4_20),.acc(r4_20),.res(r4_21),.clk(clk),.wout(w4_21));
	PE pe4_22(.x(x22),.w(w4_21),.acc(r4_21),.res(r4_22),.clk(clk),.wout(w4_22));
	PE pe4_23(.x(x23),.w(w4_22),.acc(r4_22),.res(r4_23),.clk(clk),.wout(w4_23));
	PE pe4_24(.x(x24),.w(w4_23),.acc(r4_23),.res(r4_24),.clk(clk),.wout(w4_24));
	PE pe4_25(.x(x25),.w(w4_24),.acc(r4_24),.res(r4_25),.clk(clk),.wout(w4_25));
	PE pe4_26(.x(x26),.w(w4_25),.acc(r4_25),.res(r4_26),.clk(clk),.wout(w4_26));
	PE pe4_27(.x(x27),.w(w4_26),.acc(r4_26),.res(r4_27),.clk(clk),.wout(w4_27));
	PE pe4_28(.x(x28),.w(w4_27),.acc(r4_27),.res(r4_28),.clk(clk),.wout(w4_28));
	PE pe4_29(.x(x29),.w(w4_28),.acc(r4_28),.res(r4_29),.clk(clk),.wout(w4_29));
	PE pe4_30(.x(x30),.w(w4_29),.acc(r4_29),.res(r4_30),.clk(clk),.wout(w4_30));
	PE pe4_31(.x(x31),.w(w4_30),.acc(r4_30),.res(r4_31),.clk(clk),.wout(w4_31));
	PE pe4_32(.x(x32),.w(w4_31),.acc(r4_31),.res(r4_32),.clk(clk),.wout(w4_32));
	PE pe4_33(.x(x33),.w(w4_32),.acc(r4_32),.res(r4_33),.clk(clk),.wout(w4_33));
	PE pe4_34(.x(x34),.w(w4_33),.acc(r4_33),.res(r4_34),.clk(clk),.wout(w4_34));
	PE pe4_35(.x(x35),.w(w4_34),.acc(r4_34),.res(r4_35),.clk(clk),.wout(w4_35));
	PE pe4_36(.x(x36),.w(w4_35),.acc(r4_35),.res(r4_36),.clk(clk),.wout(w4_36));
	PE pe4_37(.x(x37),.w(w4_36),.acc(r4_36),.res(r4_37),.clk(clk),.wout(w4_37));
	PE pe4_38(.x(x38),.w(w4_37),.acc(r4_37),.res(r4_38),.clk(clk),.wout(w4_38));
	PE pe4_39(.x(x39),.w(w4_38),.acc(r4_38),.res(r4_39),.clk(clk),.wout(w4_39));
	PE pe4_40(.x(x40),.w(w4_39),.acc(r4_39),.res(r4_40),.clk(clk),.wout(w4_40));
	PE pe4_41(.x(x41),.w(w4_40),.acc(r4_40),.res(r4_41),.clk(clk),.wout(w4_41));
	PE pe4_42(.x(x42),.w(w4_41),.acc(r4_41),.res(r4_42),.clk(clk),.wout(w4_42));
	PE pe4_43(.x(x43),.w(w4_42),.acc(r4_42),.res(r4_43),.clk(clk),.wout(w4_43));
	PE pe4_44(.x(x44),.w(w4_43),.acc(r4_43),.res(r4_44),.clk(clk),.wout(w4_44));
	PE pe4_45(.x(x45),.w(w4_44),.acc(r4_44),.res(r4_45),.clk(clk),.wout(w4_45));
	PE pe4_46(.x(x46),.w(w4_45),.acc(r4_45),.res(r4_46),.clk(clk),.wout(w4_46));
	PE pe4_47(.x(x47),.w(w4_46),.acc(r4_46),.res(r4_47),.clk(clk),.wout(w4_47));
	PE pe4_48(.x(x48),.w(w4_47),.acc(r4_47),.res(r4_48),.clk(clk),.wout(w4_48));
	PE pe4_49(.x(x49),.w(w4_48),.acc(r4_48),.res(r4_49),.clk(clk),.wout(w4_49));
	PE pe4_50(.x(x50),.w(w4_49),.acc(r4_49),.res(r4_50),.clk(clk),.wout(w4_50));
	PE pe4_51(.x(x51),.w(w4_50),.acc(r4_50),.res(r4_51),.clk(clk),.wout(w4_51));
	PE pe4_52(.x(x52),.w(w4_51),.acc(r4_51),.res(r4_52),.clk(clk),.wout(w4_52));
	PE pe4_53(.x(x53),.w(w4_52),.acc(r4_52),.res(r4_53),.clk(clk),.wout(w4_53));
	PE pe4_54(.x(x54),.w(w4_53),.acc(r4_53),.res(r4_54),.clk(clk),.wout(w4_54));
	PE pe4_55(.x(x55),.w(w4_54),.acc(r4_54),.res(r4_55),.clk(clk),.wout(w4_55));
	PE pe4_56(.x(x56),.w(w4_55),.acc(r4_55),.res(r4_56),.clk(clk),.wout(w4_56));
	PE pe4_57(.x(x57),.w(w4_56),.acc(r4_56),.res(r4_57),.clk(clk),.wout(w4_57));
	PE pe4_58(.x(x58),.w(w4_57),.acc(r4_57),.res(r4_58),.clk(clk),.wout(w4_58));
	PE pe4_59(.x(x59),.w(w4_58),.acc(r4_58),.res(r4_59),.clk(clk),.wout(w4_59));
	PE pe4_60(.x(x60),.w(w4_59),.acc(r4_59),.res(r4_60),.clk(clk),.wout(w4_60));
	PE pe4_61(.x(x61),.w(w4_60),.acc(r4_60),.res(r4_61),.clk(clk),.wout(w4_61));
	PE pe4_62(.x(x62),.w(w4_61),.acc(r4_61),.res(r4_62),.clk(clk),.wout(w4_62));
	PE pe4_63(.x(x63),.w(w4_62),.acc(r4_62),.res(r4_63),.clk(clk),.wout(w4_63));
	PE pe4_64(.x(x64),.w(w4_63),.acc(r4_63),.res(r4_64),.clk(clk),.wout(w4_64));
	PE pe4_65(.x(x65),.w(w4_64),.acc(r4_64),.res(r4_65),.clk(clk),.wout(w4_65));
	PE pe4_66(.x(x66),.w(w4_65),.acc(r4_65),.res(r4_66),.clk(clk),.wout(w4_66));
	PE pe4_67(.x(x67),.w(w4_66),.acc(r4_66),.res(r4_67),.clk(clk),.wout(w4_67));
	PE pe4_68(.x(x68),.w(w4_67),.acc(r4_67),.res(r4_68),.clk(clk),.wout(w4_68));
	PE pe4_69(.x(x69),.w(w4_68),.acc(r4_68),.res(r4_69),.clk(clk),.wout(w4_69));
	PE pe4_70(.x(x70),.w(w4_69),.acc(r4_69),.res(r4_70),.clk(clk),.wout(w4_70));
	PE pe4_71(.x(x71),.w(w4_70),.acc(r4_70),.res(r4_71),.clk(clk),.wout(w4_71));
	PE pe4_72(.x(x72),.w(w4_71),.acc(r4_71),.res(r4_72),.clk(clk),.wout(w4_72));
	PE pe4_73(.x(x73),.w(w4_72),.acc(r4_72),.res(r4_73),.clk(clk),.wout(w4_73));
	PE pe4_74(.x(x74),.w(w4_73),.acc(r4_73),.res(r4_74),.clk(clk),.wout(w4_74));
	PE pe4_75(.x(x75),.w(w4_74),.acc(r4_74),.res(r4_75),.clk(clk),.wout(w4_75));
	PE pe4_76(.x(x76),.w(w4_75),.acc(r4_75),.res(r4_76),.clk(clk),.wout(w4_76));
	PE pe4_77(.x(x77),.w(w4_76),.acc(r4_76),.res(r4_77),.clk(clk),.wout(w4_77));
	PE pe4_78(.x(x78),.w(w4_77),.acc(r4_77),.res(r4_78),.clk(clk),.wout(w4_78));
	PE pe4_79(.x(x79),.w(w4_78),.acc(r4_78),.res(r4_79),.clk(clk),.wout(w4_79));
	PE pe4_80(.x(x80),.w(w4_79),.acc(r4_79),.res(r4_80),.clk(clk),.wout(w4_80));
	PE pe4_81(.x(x81),.w(w4_80),.acc(r4_80),.res(r4_81),.clk(clk),.wout(w4_81));
	PE pe4_82(.x(x82),.w(w4_81),.acc(r4_81),.res(r4_82),.clk(clk),.wout(w4_82));
	PE pe4_83(.x(x83),.w(w4_82),.acc(r4_82),.res(r4_83),.clk(clk),.wout(w4_83));
	PE pe4_84(.x(x84),.w(w4_83),.acc(r4_83),.res(r4_84),.clk(clk),.wout(w4_84));
	PE pe4_85(.x(x85),.w(w4_84),.acc(r4_84),.res(r4_85),.clk(clk),.wout(w4_85));
	PE pe4_86(.x(x86),.w(w4_85),.acc(r4_85),.res(r4_86),.clk(clk),.wout(w4_86));
	PE pe4_87(.x(x87),.w(w4_86),.acc(r4_86),.res(r4_87),.clk(clk),.wout(w4_87));
	PE pe4_88(.x(x88),.w(w4_87),.acc(r4_87),.res(r4_88),.clk(clk),.wout(w4_88));
	PE pe4_89(.x(x89),.w(w4_88),.acc(r4_88),.res(r4_89),.clk(clk),.wout(w4_89));
	PE pe4_90(.x(x90),.w(w4_89),.acc(r4_89),.res(r4_90),.clk(clk),.wout(w4_90));
	PE pe4_91(.x(x91),.w(w4_90),.acc(r4_90),.res(r4_91),.clk(clk),.wout(w4_91));
	PE pe4_92(.x(x92),.w(w4_91),.acc(r4_91),.res(r4_92),.clk(clk),.wout(w4_92));
	PE pe4_93(.x(x93),.w(w4_92),.acc(r4_92),.res(r4_93),.clk(clk),.wout(w4_93));
	PE pe4_94(.x(x94),.w(w4_93),.acc(r4_93),.res(r4_94),.clk(clk),.wout(w4_94));
	PE pe4_95(.x(x95),.w(w4_94),.acc(r4_94),.res(r4_95),.clk(clk),.wout(w4_95));
	PE pe4_96(.x(x96),.w(w4_95),.acc(r4_95),.res(r4_96),.clk(clk),.wout(w4_96));
	PE pe4_97(.x(x97),.w(w4_96),.acc(r4_96),.res(r4_97),.clk(clk),.wout(w4_97));
	PE pe4_98(.x(x98),.w(w4_97),.acc(r4_97),.res(r4_98),.clk(clk),.wout(w4_98));
	PE pe4_99(.x(x99),.w(w4_98),.acc(r4_98),.res(r4_99),.clk(clk),.wout(w4_99));
	PE pe4_100(.x(x100),.w(w4_99),.acc(r4_99),.res(r4_100),.clk(clk),.wout(w4_100));
	PE pe4_101(.x(x101),.w(w4_100),.acc(r4_100),.res(r4_101),.clk(clk),.wout(w4_101));
	PE pe4_102(.x(x102),.w(w4_101),.acc(r4_101),.res(r4_102),.clk(clk),.wout(w4_102));
	PE pe4_103(.x(x103),.w(w4_102),.acc(r4_102),.res(r4_103),.clk(clk),.wout(w4_103));
	PE pe4_104(.x(x104),.w(w4_103),.acc(r4_103),.res(r4_104),.clk(clk),.wout(w4_104));
	PE pe4_105(.x(x105),.w(w4_104),.acc(r4_104),.res(r4_105),.clk(clk),.wout(w4_105));
	PE pe4_106(.x(x106),.w(w4_105),.acc(r4_105),.res(r4_106),.clk(clk),.wout(w4_106));
	PE pe4_107(.x(x107),.w(w4_106),.acc(r4_106),.res(r4_107),.clk(clk),.wout(w4_107));
	PE pe4_108(.x(x108),.w(w4_107),.acc(r4_107),.res(r4_108),.clk(clk),.wout(w4_108));
	PE pe4_109(.x(x109),.w(w4_108),.acc(r4_108),.res(r4_109),.clk(clk),.wout(w4_109));
	PE pe4_110(.x(x110),.w(w4_109),.acc(r4_109),.res(r4_110),.clk(clk),.wout(w4_110));
	PE pe4_111(.x(x111),.w(w4_110),.acc(r4_110),.res(r4_111),.clk(clk),.wout(w4_111));
	PE pe4_112(.x(x112),.w(w4_111),.acc(r4_111),.res(r4_112),.clk(clk),.wout(w4_112));
	PE pe4_113(.x(x113),.w(w4_112),.acc(r4_112),.res(r4_113),.clk(clk),.wout(w4_113));
	PE pe4_114(.x(x114),.w(w4_113),.acc(r4_113),.res(r4_114),.clk(clk),.wout(w4_114));
	PE pe4_115(.x(x115),.w(w4_114),.acc(r4_114),.res(r4_115),.clk(clk),.wout(w4_115));
	PE pe4_116(.x(x116),.w(w4_115),.acc(r4_115),.res(r4_116),.clk(clk),.wout(w4_116));
	PE pe4_117(.x(x117),.w(w4_116),.acc(r4_116),.res(r4_117),.clk(clk),.wout(w4_117));
	PE pe4_118(.x(x118),.w(w4_117),.acc(r4_117),.res(r4_118),.clk(clk),.wout(w4_118));
	PE pe4_119(.x(x119),.w(w4_118),.acc(r4_118),.res(r4_119),.clk(clk),.wout(w4_119));
	PE pe4_120(.x(x120),.w(w4_119),.acc(r4_119),.res(r4_120),.clk(clk),.wout(w4_120));
	PE pe4_121(.x(x121),.w(w4_120),.acc(r4_120),.res(r4_121),.clk(clk),.wout(w4_121));
	PE pe4_122(.x(x122),.w(w4_121),.acc(r4_121),.res(r4_122),.clk(clk),.wout(w4_122));
	PE pe4_123(.x(x123),.w(w4_122),.acc(r4_122),.res(r4_123),.clk(clk),.wout(w4_123));
	PE pe4_124(.x(x124),.w(w4_123),.acc(r4_123),.res(r4_124),.clk(clk),.wout(w4_124));
	PE pe4_125(.x(x125),.w(w4_124),.acc(r4_124),.res(r4_125),.clk(clk),.wout(w4_125));
	PE pe4_126(.x(x126),.w(w4_125),.acc(r4_125),.res(r4_126),.clk(clk),.wout(w4_126));
	PE pe4_127(.x(x127),.w(w4_126),.acc(r4_126),.res(result4),.clk(clk),.wout(weight4));

	PE pe5_0(.x(x0),.w(w5),.acc(32'h0),.res(r5_0),.clk(clk),.wout(w5_0));
	PE pe5_1(.x(x1),.w(w5_0),.acc(r5_0),.res(r5_1),.clk(clk),.wout(w5_1));
	PE pe5_2(.x(x2),.w(w5_1),.acc(r5_1),.res(r5_2),.clk(clk),.wout(w5_2));
	PE pe5_3(.x(x3),.w(w5_2),.acc(r5_2),.res(r5_3),.clk(clk),.wout(w5_3));
	PE pe5_4(.x(x4),.w(w5_3),.acc(r5_3),.res(r5_4),.clk(clk),.wout(w5_4));
	PE pe5_5(.x(x5),.w(w5_4),.acc(r5_4),.res(r5_5),.clk(clk),.wout(w5_5));
	PE pe5_6(.x(x6),.w(w5_5),.acc(r5_5),.res(r5_6),.clk(clk),.wout(w5_6));
	PE pe5_7(.x(x7),.w(w5_6),.acc(r5_6),.res(r5_7),.clk(clk),.wout(w5_7));
	PE pe5_8(.x(x8),.w(w5_7),.acc(r5_7),.res(r5_8),.clk(clk),.wout(w5_8));
	PE pe5_9(.x(x9),.w(w5_8),.acc(r5_8),.res(r5_9),.clk(clk),.wout(w5_9));
	PE pe5_10(.x(x10),.w(w5_9),.acc(r5_9),.res(r5_10),.clk(clk),.wout(w5_10));
	PE pe5_11(.x(x11),.w(w5_10),.acc(r5_10),.res(r5_11),.clk(clk),.wout(w5_11));
	PE pe5_12(.x(x12),.w(w5_11),.acc(r5_11),.res(r5_12),.clk(clk),.wout(w5_12));
	PE pe5_13(.x(x13),.w(w5_12),.acc(r5_12),.res(r5_13),.clk(clk),.wout(w5_13));
	PE pe5_14(.x(x14),.w(w5_13),.acc(r5_13),.res(r5_14),.clk(clk),.wout(w5_14));
	PE pe5_15(.x(x15),.w(w5_14),.acc(r5_14),.res(r5_15),.clk(clk),.wout(w5_15));
	PE pe5_16(.x(x16),.w(w5_15),.acc(r5_15),.res(r5_16),.clk(clk),.wout(w5_16));
	PE pe5_17(.x(x17),.w(w5_16),.acc(r5_16),.res(r5_17),.clk(clk),.wout(w5_17));
	PE pe5_18(.x(x18),.w(w5_17),.acc(r5_17),.res(r5_18),.clk(clk),.wout(w5_18));
	PE pe5_19(.x(x19),.w(w5_18),.acc(r5_18),.res(r5_19),.clk(clk),.wout(w5_19));
	PE pe5_20(.x(x20),.w(w5_19),.acc(r5_19),.res(r5_20),.clk(clk),.wout(w5_20));
	PE pe5_21(.x(x21),.w(w5_20),.acc(r5_20),.res(r5_21),.clk(clk),.wout(w5_21));
	PE pe5_22(.x(x22),.w(w5_21),.acc(r5_21),.res(r5_22),.clk(clk),.wout(w5_22));
	PE pe5_23(.x(x23),.w(w5_22),.acc(r5_22),.res(r5_23),.clk(clk),.wout(w5_23));
	PE pe5_24(.x(x24),.w(w5_23),.acc(r5_23),.res(r5_24),.clk(clk),.wout(w5_24));
	PE pe5_25(.x(x25),.w(w5_24),.acc(r5_24),.res(r5_25),.clk(clk),.wout(w5_25));
	PE pe5_26(.x(x26),.w(w5_25),.acc(r5_25),.res(r5_26),.clk(clk),.wout(w5_26));
	PE pe5_27(.x(x27),.w(w5_26),.acc(r5_26),.res(r5_27),.clk(clk),.wout(w5_27));
	PE pe5_28(.x(x28),.w(w5_27),.acc(r5_27),.res(r5_28),.clk(clk),.wout(w5_28));
	PE pe5_29(.x(x29),.w(w5_28),.acc(r5_28),.res(r5_29),.clk(clk),.wout(w5_29));
	PE pe5_30(.x(x30),.w(w5_29),.acc(r5_29),.res(r5_30),.clk(clk),.wout(w5_30));
	PE pe5_31(.x(x31),.w(w5_30),.acc(r5_30),.res(r5_31),.clk(clk),.wout(w5_31));
	PE pe5_32(.x(x32),.w(w5_31),.acc(r5_31),.res(r5_32),.clk(clk),.wout(w5_32));
	PE pe5_33(.x(x33),.w(w5_32),.acc(r5_32),.res(r5_33),.clk(clk),.wout(w5_33));
	PE pe5_34(.x(x34),.w(w5_33),.acc(r5_33),.res(r5_34),.clk(clk),.wout(w5_34));
	PE pe5_35(.x(x35),.w(w5_34),.acc(r5_34),.res(r5_35),.clk(clk),.wout(w5_35));
	PE pe5_36(.x(x36),.w(w5_35),.acc(r5_35),.res(r5_36),.clk(clk),.wout(w5_36));
	PE pe5_37(.x(x37),.w(w5_36),.acc(r5_36),.res(r5_37),.clk(clk),.wout(w5_37));
	PE pe5_38(.x(x38),.w(w5_37),.acc(r5_37),.res(r5_38),.clk(clk),.wout(w5_38));
	PE pe5_39(.x(x39),.w(w5_38),.acc(r5_38),.res(r5_39),.clk(clk),.wout(w5_39));
	PE pe5_40(.x(x40),.w(w5_39),.acc(r5_39),.res(r5_40),.clk(clk),.wout(w5_40));
	PE pe5_41(.x(x41),.w(w5_40),.acc(r5_40),.res(r5_41),.clk(clk),.wout(w5_41));
	PE pe5_42(.x(x42),.w(w5_41),.acc(r5_41),.res(r5_42),.clk(clk),.wout(w5_42));
	PE pe5_43(.x(x43),.w(w5_42),.acc(r5_42),.res(r5_43),.clk(clk),.wout(w5_43));
	PE pe5_44(.x(x44),.w(w5_43),.acc(r5_43),.res(r5_44),.clk(clk),.wout(w5_44));
	PE pe5_45(.x(x45),.w(w5_44),.acc(r5_44),.res(r5_45),.clk(clk),.wout(w5_45));
	PE pe5_46(.x(x46),.w(w5_45),.acc(r5_45),.res(r5_46),.clk(clk),.wout(w5_46));
	PE pe5_47(.x(x47),.w(w5_46),.acc(r5_46),.res(r5_47),.clk(clk),.wout(w5_47));
	PE pe5_48(.x(x48),.w(w5_47),.acc(r5_47),.res(r5_48),.clk(clk),.wout(w5_48));
	PE pe5_49(.x(x49),.w(w5_48),.acc(r5_48),.res(r5_49),.clk(clk),.wout(w5_49));
	PE pe5_50(.x(x50),.w(w5_49),.acc(r5_49),.res(r5_50),.clk(clk),.wout(w5_50));
	PE pe5_51(.x(x51),.w(w5_50),.acc(r5_50),.res(r5_51),.clk(clk),.wout(w5_51));
	PE pe5_52(.x(x52),.w(w5_51),.acc(r5_51),.res(r5_52),.clk(clk),.wout(w5_52));
	PE pe5_53(.x(x53),.w(w5_52),.acc(r5_52),.res(r5_53),.clk(clk),.wout(w5_53));
	PE pe5_54(.x(x54),.w(w5_53),.acc(r5_53),.res(r5_54),.clk(clk),.wout(w5_54));
	PE pe5_55(.x(x55),.w(w5_54),.acc(r5_54),.res(r5_55),.clk(clk),.wout(w5_55));
	PE pe5_56(.x(x56),.w(w5_55),.acc(r5_55),.res(r5_56),.clk(clk),.wout(w5_56));
	PE pe5_57(.x(x57),.w(w5_56),.acc(r5_56),.res(r5_57),.clk(clk),.wout(w5_57));
	PE pe5_58(.x(x58),.w(w5_57),.acc(r5_57),.res(r5_58),.clk(clk),.wout(w5_58));
	PE pe5_59(.x(x59),.w(w5_58),.acc(r5_58),.res(r5_59),.clk(clk),.wout(w5_59));
	PE pe5_60(.x(x60),.w(w5_59),.acc(r5_59),.res(r5_60),.clk(clk),.wout(w5_60));
	PE pe5_61(.x(x61),.w(w5_60),.acc(r5_60),.res(r5_61),.clk(clk),.wout(w5_61));
	PE pe5_62(.x(x62),.w(w5_61),.acc(r5_61),.res(r5_62),.clk(clk),.wout(w5_62));
	PE pe5_63(.x(x63),.w(w5_62),.acc(r5_62),.res(r5_63),.clk(clk),.wout(w5_63));
	PE pe5_64(.x(x64),.w(w5_63),.acc(r5_63),.res(r5_64),.clk(clk),.wout(w5_64));
	PE pe5_65(.x(x65),.w(w5_64),.acc(r5_64),.res(r5_65),.clk(clk),.wout(w5_65));
	PE pe5_66(.x(x66),.w(w5_65),.acc(r5_65),.res(r5_66),.clk(clk),.wout(w5_66));
	PE pe5_67(.x(x67),.w(w5_66),.acc(r5_66),.res(r5_67),.clk(clk),.wout(w5_67));
	PE pe5_68(.x(x68),.w(w5_67),.acc(r5_67),.res(r5_68),.clk(clk),.wout(w5_68));
	PE pe5_69(.x(x69),.w(w5_68),.acc(r5_68),.res(r5_69),.clk(clk),.wout(w5_69));
	PE pe5_70(.x(x70),.w(w5_69),.acc(r5_69),.res(r5_70),.clk(clk),.wout(w5_70));
	PE pe5_71(.x(x71),.w(w5_70),.acc(r5_70),.res(r5_71),.clk(clk),.wout(w5_71));
	PE pe5_72(.x(x72),.w(w5_71),.acc(r5_71),.res(r5_72),.clk(clk),.wout(w5_72));
	PE pe5_73(.x(x73),.w(w5_72),.acc(r5_72),.res(r5_73),.clk(clk),.wout(w5_73));
	PE pe5_74(.x(x74),.w(w5_73),.acc(r5_73),.res(r5_74),.clk(clk),.wout(w5_74));
	PE pe5_75(.x(x75),.w(w5_74),.acc(r5_74),.res(r5_75),.clk(clk),.wout(w5_75));
	PE pe5_76(.x(x76),.w(w5_75),.acc(r5_75),.res(r5_76),.clk(clk),.wout(w5_76));
	PE pe5_77(.x(x77),.w(w5_76),.acc(r5_76),.res(r5_77),.clk(clk),.wout(w5_77));
	PE pe5_78(.x(x78),.w(w5_77),.acc(r5_77),.res(r5_78),.clk(clk),.wout(w5_78));
	PE pe5_79(.x(x79),.w(w5_78),.acc(r5_78),.res(r5_79),.clk(clk),.wout(w5_79));
	PE pe5_80(.x(x80),.w(w5_79),.acc(r5_79),.res(r5_80),.clk(clk),.wout(w5_80));
	PE pe5_81(.x(x81),.w(w5_80),.acc(r5_80),.res(r5_81),.clk(clk),.wout(w5_81));
	PE pe5_82(.x(x82),.w(w5_81),.acc(r5_81),.res(r5_82),.clk(clk),.wout(w5_82));
	PE pe5_83(.x(x83),.w(w5_82),.acc(r5_82),.res(r5_83),.clk(clk),.wout(w5_83));
	PE pe5_84(.x(x84),.w(w5_83),.acc(r5_83),.res(r5_84),.clk(clk),.wout(w5_84));
	PE pe5_85(.x(x85),.w(w5_84),.acc(r5_84),.res(r5_85),.clk(clk),.wout(w5_85));
	PE pe5_86(.x(x86),.w(w5_85),.acc(r5_85),.res(r5_86),.clk(clk),.wout(w5_86));
	PE pe5_87(.x(x87),.w(w5_86),.acc(r5_86),.res(r5_87),.clk(clk),.wout(w5_87));
	PE pe5_88(.x(x88),.w(w5_87),.acc(r5_87),.res(r5_88),.clk(clk),.wout(w5_88));
	PE pe5_89(.x(x89),.w(w5_88),.acc(r5_88),.res(r5_89),.clk(clk),.wout(w5_89));
	PE pe5_90(.x(x90),.w(w5_89),.acc(r5_89),.res(r5_90),.clk(clk),.wout(w5_90));
	PE pe5_91(.x(x91),.w(w5_90),.acc(r5_90),.res(r5_91),.clk(clk),.wout(w5_91));
	PE pe5_92(.x(x92),.w(w5_91),.acc(r5_91),.res(r5_92),.clk(clk),.wout(w5_92));
	PE pe5_93(.x(x93),.w(w5_92),.acc(r5_92),.res(r5_93),.clk(clk),.wout(w5_93));
	PE pe5_94(.x(x94),.w(w5_93),.acc(r5_93),.res(r5_94),.clk(clk),.wout(w5_94));
	PE pe5_95(.x(x95),.w(w5_94),.acc(r5_94),.res(r5_95),.clk(clk),.wout(w5_95));
	PE pe5_96(.x(x96),.w(w5_95),.acc(r5_95),.res(r5_96),.clk(clk),.wout(w5_96));
	PE pe5_97(.x(x97),.w(w5_96),.acc(r5_96),.res(r5_97),.clk(clk),.wout(w5_97));
	PE pe5_98(.x(x98),.w(w5_97),.acc(r5_97),.res(r5_98),.clk(clk),.wout(w5_98));
	PE pe5_99(.x(x99),.w(w5_98),.acc(r5_98),.res(r5_99),.clk(clk),.wout(w5_99));
	PE pe5_100(.x(x100),.w(w5_99),.acc(r5_99),.res(r5_100),.clk(clk),.wout(w5_100));
	PE pe5_101(.x(x101),.w(w5_100),.acc(r5_100),.res(r5_101),.clk(clk),.wout(w5_101));
	PE pe5_102(.x(x102),.w(w5_101),.acc(r5_101),.res(r5_102),.clk(clk),.wout(w5_102));
	PE pe5_103(.x(x103),.w(w5_102),.acc(r5_102),.res(r5_103),.clk(clk),.wout(w5_103));
	PE pe5_104(.x(x104),.w(w5_103),.acc(r5_103),.res(r5_104),.clk(clk),.wout(w5_104));
	PE pe5_105(.x(x105),.w(w5_104),.acc(r5_104),.res(r5_105),.clk(clk),.wout(w5_105));
	PE pe5_106(.x(x106),.w(w5_105),.acc(r5_105),.res(r5_106),.clk(clk),.wout(w5_106));
	PE pe5_107(.x(x107),.w(w5_106),.acc(r5_106),.res(r5_107),.clk(clk),.wout(w5_107));
	PE pe5_108(.x(x108),.w(w5_107),.acc(r5_107),.res(r5_108),.clk(clk),.wout(w5_108));
	PE pe5_109(.x(x109),.w(w5_108),.acc(r5_108),.res(r5_109),.clk(clk),.wout(w5_109));
	PE pe5_110(.x(x110),.w(w5_109),.acc(r5_109),.res(r5_110),.clk(clk),.wout(w5_110));
	PE pe5_111(.x(x111),.w(w5_110),.acc(r5_110),.res(r5_111),.clk(clk),.wout(w5_111));
	PE pe5_112(.x(x112),.w(w5_111),.acc(r5_111),.res(r5_112),.clk(clk),.wout(w5_112));
	PE pe5_113(.x(x113),.w(w5_112),.acc(r5_112),.res(r5_113),.clk(clk),.wout(w5_113));
	PE pe5_114(.x(x114),.w(w5_113),.acc(r5_113),.res(r5_114),.clk(clk),.wout(w5_114));
	PE pe5_115(.x(x115),.w(w5_114),.acc(r5_114),.res(r5_115),.clk(clk),.wout(w5_115));
	PE pe5_116(.x(x116),.w(w5_115),.acc(r5_115),.res(r5_116),.clk(clk),.wout(w5_116));
	PE pe5_117(.x(x117),.w(w5_116),.acc(r5_116),.res(r5_117),.clk(clk),.wout(w5_117));
	PE pe5_118(.x(x118),.w(w5_117),.acc(r5_117),.res(r5_118),.clk(clk),.wout(w5_118));
	PE pe5_119(.x(x119),.w(w5_118),.acc(r5_118),.res(r5_119),.clk(clk),.wout(w5_119));
	PE pe5_120(.x(x120),.w(w5_119),.acc(r5_119),.res(r5_120),.clk(clk),.wout(w5_120));
	PE pe5_121(.x(x121),.w(w5_120),.acc(r5_120),.res(r5_121),.clk(clk),.wout(w5_121));
	PE pe5_122(.x(x122),.w(w5_121),.acc(r5_121),.res(r5_122),.clk(clk),.wout(w5_122));
	PE pe5_123(.x(x123),.w(w5_122),.acc(r5_122),.res(r5_123),.clk(clk),.wout(w5_123));
	PE pe5_124(.x(x124),.w(w5_123),.acc(r5_123),.res(r5_124),.clk(clk),.wout(w5_124));
	PE pe5_125(.x(x125),.w(w5_124),.acc(r5_124),.res(r5_125),.clk(clk),.wout(w5_125));
	PE pe5_126(.x(x126),.w(w5_125),.acc(r5_125),.res(r5_126),.clk(clk),.wout(w5_126));
	PE pe5_127(.x(x127),.w(w5_126),.acc(r5_126),.res(result5),.clk(clk),.wout(weight5));

	PE pe6_0(.x(x0),.w(w6),.acc(32'h0),.res(r6_0),.clk(clk),.wout(w6_0));
	PE pe6_1(.x(x1),.w(w6_0),.acc(r6_0),.res(r6_1),.clk(clk),.wout(w6_1));
	PE pe6_2(.x(x2),.w(w6_1),.acc(r6_1),.res(r6_2),.clk(clk),.wout(w6_2));
	PE pe6_3(.x(x3),.w(w6_2),.acc(r6_2),.res(r6_3),.clk(clk),.wout(w6_3));
	PE pe6_4(.x(x4),.w(w6_3),.acc(r6_3),.res(r6_4),.clk(clk),.wout(w6_4));
	PE pe6_5(.x(x5),.w(w6_4),.acc(r6_4),.res(r6_5),.clk(clk),.wout(w6_5));
	PE pe6_6(.x(x6),.w(w6_5),.acc(r6_5),.res(r6_6),.clk(clk),.wout(w6_6));
	PE pe6_7(.x(x7),.w(w6_6),.acc(r6_6),.res(r6_7),.clk(clk),.wout(w6_7));
	PE pe6_8(.x(x8),.w(w6_7),.acc(r6_7),.res(r6_8),.clk(clk),.wout(w6_8));
	PE pe6_9(.x(x9),.w(w6_8),.acc(r6_8),.res(r6_9),.clk(clk),.wout(w6_9));
	PE pe6_10(.x(x10),.w(w6_9),.acc(r6_9),.res(r6_10),.clk(clk),.wout(w6_10));
	PE pe6_11(.x(x11),.w(w6_10),.acc(r6_10),.res(r6_11),.clk(clk),.wout(w6_11));
	PE pe6_12(.x(x12),.w(w6_11),.acc(r6_11),.res(r6_12),.clk(clk),.wout(w6_12));
	PE pe6_13(.x(x13),.w(w6_12),.acc(r6_12),.res(r6_13),.clk(clk),.wout(w6_13));
	PE pe6_14(.x(x14),.w(w6_13),.acc(r6_13),.res(r6_14),.clk(clk),.wout(w6_14));
	PE pe6_15(.x(x15),.w(w6_14),.acc(r6_14),.res(r6_15),.clk(clk),.wout(w6_15));
	PE pe6_16(.x(x16),.w(w6_15),.acc(r6_15),.res(r6_16),.clk(clk),.wout(w6_16));
	PE pe6_17(.x(x17),.w(w6_16),.acc(r6_16),.res(r6_17),.clk(clk),.wout(w6_17));
	PE pe6_18(.x(x18),.w(w6_17),.acc(r6_17),.res(r6_18),.clk(clk),.wout(w6_18));
	PE pe6_19(.x(x19),.w(w6_18),.acc(r6_18),.res(r6_19),.clk(clk),.wout(w6_19));
	PE pe6_20(.x(x20),.w(w6_19),.acc(r6_19),.res(r6_20),.clk(clk),.wout(w6_20));
	PE pe6_21(.x(x21),.w(w6_20),.acc(r6_20),.res(r6_21),.clk(clk),.wout(w6_21));
	PE pe6_22(.x(x22),.w(w6_21),.acc(r6_21),.res(r6_22),.clk(clk),.wout(w6_22));
	PE pe6_23(.x(x23),.w(w6_22),.acc(r6_22),.res(r6_23),.clk(clk),.wout(w6_23));
	PE pe6_24(.x(x24),.w(w6_23),.acc(r6_23),.res(r6_24),.clk(clk),.wout(w6_24));
	PE pe6_25(.x(x25),.w(w6_24),.acc(r6_24),.res(r6_25),.clk(clk),.wout(w6_25));
	PE pe6_26(.x(x26),.w(w6_25),.acc(r6_25),.res(r6_26),.clk(clk),.wout(w6_26));
	PE pe6_27(.x(x27),.w(w6_26),.acc(r6_26),.res(r6_27),.clk(clk),.wout(w6_27));
	PE pe6_28(.x(x28),.w(w6_27),.acc(r6_27),.res(r6_28),.clk(clk),.wout(w6_28));
	PE pe6_29(.x(x29),.w(w6_28),.acc(r6_28),.res(r6_29),.clk(clk),.wout(w6_29));
	PE pe6_30(.x(x30),.w(w6_29),.acc(r6_29),.res(r6_30),.clk(clk),.wout(w6_30));
	PE pe6_31(.x(x31),.w(w6_30),.acc(r6_30),.res(r6_31),.clk(clk),.wout(w6_31));
	PE pe6_32(.x(x32),.w(w6_31),.acc(r6_31),.res(r6_32),.clk(clk),.wout(w6_32));
	PE pe6_33(.x(x33),.w(w6_32),.acc(r6_32),.res(r6_33),.clk(clk),.wout(w6_33));
	PE pe6_34(.x(x34),.w(w6_33),.acc(r6_33),.res(r6_34),.clk(clk),.wout(w6_34));
	PE pe6_35(.x(x35),.w(w6_34),.acc(r6_34),.res(r6_35),.clk(clk),.wout(w6_35));
	PE pe6_36(.x(x36),.w(w6_35),.acc(r6_35),.res(r6_36),.clk(clk),.wout(w6_36));
	PE pe6_37(.x(x37),.w(w6_36),.acc(r6_36),.res(r6_37),.clk(clk),.wout(w6_37));
	PE pe6_38(.x(x38),.w(w6_37),.acc(r6_37),.res(r6_38),.clk(clk),.wout(w6_38));
	PE pe6_39(.x(x39),.w(w6_38),.acc(r6_38),.res(r6_39),.clk(clk),.wout(w6_39));
	PE pe6_40(.x(x40),.w(w6_39),.acc(r6_39),.res(r6_40),.clk(clk),.wout(w6_40));
	PE pe6_41(.x(x41),.w(w6_40),.acc(r6_40),.res(r6_41),.clk(clk),.wout(w6_41));
	PE pe6_42(.x(x42),.w(w6_41),.acc(r6_41),.res(r6_42),.clk(clk),.wout(w6_42));
	PE pe6_43(.x(x43),.w(w6_42),.acc(r6_42),.res(r6_43),.clk(clk),.wout(w6_43));
	PE pe6_44(.x(x44),.w(w6_43),.acc(r6_43),.res(r6_44),.clk(clk),.wout(w6_44));
	PE pe6_45(.x(x45),.w(w6_44),.acc(r6_44),.res(r6_45),.clk(clk),.wout(w6_45));
	PE pe6_46(.x(x46),.w(w6_45),.acc(r6_45),.res(r6_46),.clk(clk),.wout(w6_46));
	PE pe6_47(.x(x47),.w(w6_46),.acc(r6_46),.res(r6_47),.clk(clk),.wout(w6_47));
	PE pe6_48(.x(x48),.w(w6_47),.acc(r6_47),.res(r6_48),.clk(clk),.wout(w6_48));
	PE pe6_49(.x(x49),.w(w6_48),.acc(r6_48),.res(r6_49),.clk(clk),.wout(w6_49));
	PE pe6_50(.x(x50),.w(w6_49),.acc(r6_49),.res(r6_50),.clk(clk),.wout(w6_50));
	PE pe6_51(.x(x51),.w(w6_50),.acc(r6_50),.res(r6_51),.clk(clk),.wout(w6_51));
	PE pe6_52(.x(x52),.w(w6_51),.acc(r6_51),.res(r6_52),.clk(clk),.wout(w6_52));
	PE pe6_53(.x(x53),.w(w6_52),.acc(r6_52),.res(r6_53),.clk(clk),.wout(w6_53));
	PE pe6_54(.x(x54),.w(w6_53),.acc(r6_53),.res(r6_54),.clk(clk),.wout(w6_54));
	PE pe6_55(.x(x55),.w(w6_54),.acc(r6_54),.res(r6_55),.clk(clk),.wout(w6_55));
	PE pe6_56(.x(x56),.w(w6_55),.acc(r6_55),.res(r6_56),.clk(clk),.wout(w6_56));
	PE pe6_57(.x(x57),.w(w6_56),.acc(r6_56),.res(r6_57),.clk(clk),.wout(w6_57));
	PE pe6_58(.x(x58),.w(w6_57),.acc(r6_57),.res(r6_58),.clk(clk),.wout(w6_58));
	PE pe6_59(.x(x59),.w(w6_58),.acc(r6_58),.res(r6_59),.clk(clk),.wout(w6_59));
	PE pe6_60(.x(x60),.w(w6_59),.acc(r6_59),.res(r6_60),.clk(clk),.wout(w6_60));
	PE pe6_61(.x(x61),.w(w6_60),.acc(r6_60),.res(r6_61),.clk(clk),.wout(w6_61));
	PE pe6_62(.x(x62),.w(w6_61),.acc(r6_61),.res(r6_62),.clk(clk),.wout(w6_62));
	PE pe6_63(.x(x63),.w(w6_62),.acc(r6_62),.res(r6_63),.clk(clk),.wout(w6_63));
	PE pe6_64(.x(x64),.w(w6_63),.acc(r6_63),.res(r6_64),.clk(clk),.wout(w6_64));
	PE pe6_65(.x(x65),.w(w6_64),.acc(r6_64),.res(r6_65),.clk(clk),.wout(w6_65));
	PE pe6_66(.x(x66),.w(w6_65),.acc(r6_65),.res(r6_66),.clk(clk),.wout(w6_66));
	PE pe6_67(.x(x67),.w(w6_66),.acc(r6_66),.res(r6_67),.clk(clk),.wout(w6_67));
	PE pe6_68(.x(x68),.w(w6_67),.acc(r6_67),.res(r6_68),.clk(clk),.wout(w6_68));
	PE pe6_69(.x(x69),.w(w6_68),.acc(r6_68),.res(r6_69),.clk(clk),.wout(w6_69));
	PE pe6_70(.x(x70),.w(w6_69),.acc(r6_69),.res(r6_70),.clk(clk),.wout(w6_70));
	PE pe6_71(.x(x71),.w(w6_70),.acc(r6_70),.res(r6_71),.clk(clk),.wout(w6_71));
	PE pe6_72(.x(x72),.w(w6_71),.acc(r6_71),.res(r6_72),.clk(clk),.wout(w6_72));
	PE pe6_73(.x(x73),.w(w6_72),.acc(r6_72),.res(r6_73),.clk(clk),.wout(w6_73));
	PE pe6_74(.x(x74),.w(w6_73),.acc(r6_73),.res(r6_74),.clk(clk),.wout(w6_74));
	PE pe6_75(.x(x75),.w(w6_74),.acc(r6_74),.res(r6_75),.clk(clk),.wout(w6_75));
	PE pe6_76(.x(x76),.w(w6_75),.acc(r6_75),.res(r6_76),.clk(clk),.wout(w6_76));
	PE pe6_77(.x(x77),.w(w6_76),.acc(r6_76),.res(r6_77),.clk(clk),.wout(w6_77));
	PE pe6_78(.x(x78),.w(w6_77),.acc(r6_77),.res(r6_78),.clk(clk),.wout(w6_78));
	PE pe6_79(.x(x79),.w(w6_78),.acc(r6_78),.res(r6_79),.clk(clk),.wout(w6_79));
	PE pe6_80(.x(x80),.w(w6_79),.acc(r6_79),.res(r6_80),.clk(clk),.wout(w6_80));
	PE pe6_81(.x(x81),.w(w6_80),.acc(r6_80),.res(r6_81),.clk(clk),.wout(w6_81));
	PE pe6_82(.x(x82),.w(w6_81),.acc(r6_81),.res(r6_82),.clk(clk),.wout(w6_82));
	PE pe6_83(.x(x83),.w(w6_82),.acc(r6_82),.res(r6_83),.clk(clk),.wout(w6_83));
	PE pe6_84(.x(x84),.w(w6_83),.acc(r6_83),.res(r6_84),.clk(clk),.wout(w6_84));
	PE pe6_85(.x(x85),.w(w6_84),.acc(r6_84),.res(r6_85),.clk(clk),.wout(w6_85));
	PE pe6_86(.x(x86),.w(w6_85),.acc(r6_85),.res(r6_86),.clk(clk),.wout(w6_86));
	PE pe6_87(.x(x87),.w(w6_86),.acc(r6_86),.res(r6_87),.clk(clk),.wout(w6_87));
	PE pe6_88(.x(x88),.w(w6_87),.acc(r6_87),.res(r6_88),.clk(clk),.wout(w6_88));
	PE pe6_89(.x(x89),.w(w6_88),.acc(r6_88),.res(r6_89),.clk(clk),.wout(w6_89));
	PE pe6_90(.x(x90),.w(w6_89),.acc(r6_89),.res(r6_90),.clk(clk),.wout(w6_90));
	PE pe6_91(.x(x91),.w(w6_90),.acc(r6_90),.res(r6_91),.clk(clk),.wout(w6_91));
	PE pe6_92(.x(x92),.w(w6_91),.acc(r6_91),.res(r6_92),.clk(clk),.wout(w6_92));
	PE pe6_93(.x(x93),.w(w6_92),.acc(r6_92),.res(r6_93),.clk(clk),.wout(w6_93));
	PE pe6_94(.x(x94),.w(w6_93),.acc(r6_93),.res(r6_94),.clk(clk),.wout(w6_94));
	PE pe6_95(.x(x95),.w(w6_94),.acc(r6_94),.res(r6_95),.clk(clk),.wout(w6_95));
	PE pe6_96(.x(x96),.w(w6_95),.acc(r6_95),.res(r6_96),.clk(clk),.wout(w6_96));
	PE pe6_97(.x(x97),.w(w6_96),.acc(r6_96),.res(r6_97),.clk(clk),.wout(w6_97));
	PE pe6_98(.x(x98),.w(w6_97),.acc(r6_97),.res(r6_98),.clk(clk),.wout(w6_98));
	PE pe6_99(.x(x99),.w(w6_98),.acc(r6_98),.res(r6_99),.clk(clk),.wout(w6_99));
	PE pe6_100(.x(x100),.w(w6_99),.acc(r6_99),.res(r6_100),.clk(clk),.wout(w6_100));
	PE pe6_101(.x(x101),.w(w6_100),.acc(r6_100),.res(r6_101),.clk(clk),.wout(w6_101));
	PE pe6_102(.x(x102),.w(w6_101),.acc(r6_101),.res(r6_102),.clk(clk),.wout(w6_102));
	PE pe6_103(.x(x103),.w(w6_102),.acc(r6_102),.res(r6_103),.clk(clk),.wout(w6_103));
	PE pe6_104(.x(x104),.w(w6_103),.acc(r6_103),.res(r6_104),.clk(clk),.wout(w6_104));
	PE pe6_105(.x(x105),.w(w6_104),.acc(r6_104),.res(r6_105),.clk(clk),.wout(w6_105));
	PE pe6_106(.x(x106),.w(w6_105),.acc(r6_105),.res(r6_106),.clk(clk),.wout(w6_106));
	PE pe6_107(.x(x107),.w(w6_106),.acc(r6_106),.res(r6_107),.clk(clk),.wout(w6_107));
	PE pe6_108(.x(x108),.w(w6_107),.acc(r6_107),.res(r6_108),.clk(clk),.wout(w6_108));
	PE pe6_109(.x(x109),.w(w6_108),.acc(r6_108),.res(r6_109),.clk(clk),.wout(w6_109));
	PE pe6_110(.x(x110),.w(w6_109),.acc(r6_109),.res(r6_110),.clk(clk),.wout(w6_110));
	PE pe6_111(.x(x111),.w(w6_110),.acc(r6_110),.res(r6_111),.clk(clk),.wout(w6_111));
	PE pe6_112(.x(x112),.w(w6_111),.acc(r6_111),.res(r6_112),.clk(clk),.wout(w6_112));
	PE pe6_113(.x(x113),.w(w6_112),.acc(r6_112),.res(r6_113),.clk(clk),.wout(w6_113));
	PE pe6_114(.x(x114),.w(w6_113),.acc(r6_113),.res(r6_114),.clk(clk),.wout(w6_114));
	PE pe6_115(.x(x115),.w(w6_114),.acc(r6_114),.res(r6_115),.clk(clk),.wout(w6_115));
	PE pe6_116(.x(x116),.w(w6_115),.acc(r6_115),.res(r6_116),.clk(clk),.wout(w6_116));
	PE pe6_117(.x(x117),.w(w6_116),.acc(r6_116),.res(r6_117),.clk(clk),.wout(w6_117));
	PE pe6_118(.x(x118),.w(w6_117),.acc(r6_117),.res(r6_118),.clk(clk),.wout(w6_118));
	PE pe6_119(.x(x119),.w(w6_118),.acc(r6_118),.res(r6_119),.clk(clk),.wout(w6_119));
	PE pe6_120(.x(x120),.w(w6_119),.acc(r6_119),.res(r6_120),.clk(clk),.wout(w6_120));
	PE pe6_121(.x(x121),.w(w6_120),.acc(r6_120),.res(r6_121),.clk(clk),.wout(w6_121));
	PE pe6_122(.x(x122),.w(w6_121),.acc(r6_121),.res(r6_122),.clk(clk),.wout(w6_122));
	PE pe6_123(.x(x123),.w(w6_122),.acc(r6_122),.res(r6_123),.clk(clk),.wout(w6_123));
	PE pe6_124(.x(x124),.w(w6_123),.acc(r6_123),.res(r6_124),.clk(clk),.wout(w6_124));
	PE pe6_125(.x(x125),.w(w6_124),.acc(r6_124),.res(r6_125),.clk(clk),.wout(w6_125));
	PE pe6_126(.x(x126),.w(w6_125),.acc(r6_125),.res(r6_126),.clk(clk),.wout(w6_126));
	PE pe6_127(.x(x127),.w(w6_126),.acc(r6_126),.res(result6),.clk(clk),.wout(weight6));

	PE pe7_0(.x(x0),.w(w7),.acc(32'h0),.res(r7_0),.clk(clk),.wout(w7_0));
	PE pe7_1(.x(x1),.w(w7_0),.acc(r7_0),.res(r7_1),.clk(clk),.wout(w7_1));
	PE pe7_2(.x(x2),.w(w7_1),.acc(r7_1),.res(r7_2),.clk(clk),.wout(w7_2));
	PE pe7_3(.x(x3),.w(w7_2),.acc(r7_2),.res(r7_3),.clk(clk),.wout(w7_3));
	PE pe7_4(.x(x4),.w(w7_3),.acc(r7_3),.res(r7_4),.clk(clk),.wout(w7_4));
	PE pe7_5(.x(x5),.w(w7_4),.acc(r7_4),.res(r7_5),.clk(clk),.wout(w7_5));
	PE pe7_6(.x(x6),.w(w7_5),.acc(r7_5),.res(r7_6),.clk(clk),.wout(w7_6));
	PE pe7_7(.x(x7),.w(w7_6),.acc(r7_6),.res(r7_7),.clk(clk),.wout(w7_7));
	PE pe7_8(.x(x8),.w(w7_7),.acc(r7_7),.res(r7_8),.clk(clk),.wout(w7_8));
	PE pe7_9(.x(x9),.w(w7_8),.acc(r7_8),.res(r7_9),.clk(clk),.wout(w7_9));
	PE pe7_10(.x(x10),.w(w7_9),.acc(r7_9),.res(r7_10),.clk(clk),.wout(w7_10));
	PE pe7_11(.x(x11),.w(w7_10),.acc(r7_10),.res(r7_11),.clk(clk),.wout(w7_11));
	PE pe7_12(.x(x12),.w(w7_11),.acc(r7_11),.res(r7_12),.clk(clk),.wout(w7_12));
	PE pe7_13(.x(x13),.w(w7_12),.acc(r7_12),.res(r7_13),.clk(clk),.wout(w7_13));
	PE pe7_14(.x(x14),.w(w7_13),.acc(r7_13),.res(r7_14),.clk(clk),.wout(w7_14));
	PE pe7_15(.x(x15),.w(w7_14),.acc(r7_14),.res(r7_15),.clk(clk),.wout(w7_15));
	PE pe7_16(.x(x16),.w(w7_15),.acc(r7_15),.res(r7_16),.clk(clk),.wout(w7_16));
	PE pe7_17(.x(x17),.w(w7_16),.acc(r7_16),.res(r7_17),.clk(clk),.wout(w7_17));
	PE pe7_18(.x(x18),.w(w7_17),.acc(r7_17),.res(r7_18),.clk(clk),.wout(w7_18));
	PE pe7_19(.x(x19),.w(w7_18),.acc(r7_18),.res(r7_19),.clk(clk),.wout(w7_19));
	PE pe7_20(.x(x20),.w(w7_19),.acc(r7_19),.res(r7_20),.clk(clk),.wout(w7_20));
	PE pe7_21(.x(x21),.w(w7_20),.acc(r7_20),.res(r7_21),.clk(clk),.wout(w7_21));
	PE pe7_22(.x(x22),.w(w7_21),.acc(r7_21),.res(r7_22),.clk(clk),.wout(w7_22));
	PE pe7_23(.x(x23),.w(w7_22),.acc(r7_22),.res(r7_23),.clk(clk),.wout(w7_23));
	PE pe7_24(.x(x24),.w(w7_23),.acc(r7_23),.res(r7_24),.clk(clk),.wout(w7_24));
	PE pe7_25(.x(x25),.w(w7_24),.acc(r7_24),.res(r7_25),.clk(clk),.wout(w7_25));
	PE pe7_26(.x(x26),.w(w7_25),.acc(r7_25),.res(r7_26),.clk(clk),.wout(w7_26));
	PE pe7_27(.x(x27),.w(w7_26),.acc(r7_26),.res(r7_27),.clk(clk),.wout(w7_27));
	PE pe7_28(.x(x28),.w(w7_27),.acc(r7_27),.res(r7_28),.clk(clk),.wout(w7_28));
	PE pe7_29(.x(x29),.w(w7_28),.acc(r7_28),.res(r7_29),.clk(clk),.wout(w7_29));
	PE pe7_30(.x(x30),.w(w7_29),.acc(r7_29),.res(r7_30),.clk(clk),.wout(w7_30));
	PE pe7_31(.x(x31),.w(w7_30),.acc(r7_30),.res(r7_31),.clk(clk),.wout(w7_31));
	PE pe7_32(.x(x32),.w(w7_31),.acc(r7_31),.res(r7_32),.clk(clk),.wout(w7_32));
	PE pe7_33(.x(x33),.w(w7_32),.acc(r7_32),.res(r7_33),.clk(clk),.wout(w7_33));
	PE pe7_34(.x(x34),.w(w7_33),.acc(r7_33),.res(r7_34),.clk(clk),.wout(w7_34));
	PE pe7_35(.x(x35),.w(w7_34),.acc(r7_34),.res(r7_35),.clk(clk),.wout(w7_35));
	PE pe7_36(.x(x36),.w(w7_35),.acc(r7_35),.res(r7_36),.clk(clk),.wout(w7_36));
	PE pe7_37(.x(x37),.w(w7_36),.acc(r7_36),.res(r7_37),.clk(clk),.wout(w7_37));
	PE pe7_38(.x(x38),.w(w7_37),.acc(r7_37),.res(r7_38),.clk(clk),.wout(w7_38));
	PE pe7_39(.x(x39),.w(w7_38),.acc(r7_38),.res(r7_39),.clk(clk),.wout(w7_39));
	PE pe7_40(.x(x40),.w(w7_39),.acc(r7_39),.res(r7_40),.clk(clk),.wout(w7_40));
	PE pe7_41(.x(x41),.w(w7_40),.acc(r7_40),.res(r7_41),.clk(clk),.wout(w7_41));
	PE pe7_42(.x(x42),.w(w7_41),.acc(r7_41),.res(r7_42),.clk(clk),.wout(w7_42));
	PE pe7_43(.x(x43),.w(w7_42),.acc(r7_42),.res(r7_43),.clk(clk),.wout(w7_43));
	PE pe7_44(.x(x44),.w(w7_43),.acc(r7_43),.res(r7_44),.clk(clk),.wout(w7_44));
	PE pe7_45(.x(x45),.w(w7_44),.acc(r7_44),.res(r7_45),.clk(clk),.wout(w7_45));
	PE pe7_46(.x(x46),.w(w7_45),.acc(r7_45),.res(r7_46),.clk(clk),.wout(w7_46));
	PE pe7_47(.x(x47),.w(w7_46),.acc(r7_46),.res(r7_47),.clk(clk),.wout(w7_47));
	PE pe7_48(.x(x48),.w(w7_47),.acc(r7_47),.res(r7_48),.clk(clk),.wout(w7_48));
	PE pe7_49(.x(x49),.w(w7_48),.acc(r7_48),.res(r7_49),.clk(clk),.wout(w7_49));
	PE pe7_50(.x(x50),.w(w7_49),.acc(r7_49),.res(r7_50),.clk(clk),.wout(w7_50));
	PE pe7_51(.x(x51),.w(w7_50),.acc(r7_50),.res(r7_51),.clk(clk),.wout(w7_51));
	PE pe7_52(.x(x52),.w(w7_51),.acc(r7_51),.res(r7_52),.clk(clk),.wout(w7_52));
	PE pe7_53(.x(x53),.w(w7_52),.acc(r7_52),.res(r7_53),.clk(clk),.wout(w7_53));
	PE pe7_54(.x(x54),.w(w7_53),.acc(r7_53),.res(r7_54),.clk(clk),.wout(w7_54));
	PE pe7_55(.x(x55),.w(w7_54),.acc(r7_54),.res(r7_55),.clk(clk),.wout(w7_55));
	PE pe7_56(.x(x56),.w(w7_55),.acc(r7_55),.res(r7_56),.clk(clk),.wout(w7_56));
	PE pe7_57(.x(x57),.w(w7_56),.acc(r7_56),.res(r7_57),.clk(clk),.wout(w7_57));
	PE pe7_58(.x(x58),.w(w7_57),.acc(r7_57),.res(r7_58),.clk(clk),.wout(w7_58));
	PE pe7_59(.x(x59),.w(w7_58),.acc(r7_58),.res(r7_59),.clk(clk),.wout(w7_59));
	PE pe7_60(.x(x60),.w(w7_59),.acc(r7_59),.res(r7_60),.clk(clk),.wout(w7_60));
	PE pe7_61(.x(x61),.w(w7_60),.acc(r7_60),.res(r7_61),.clk(clk),.wout(w7_61));
	PE pe7_62(.x(x62),.w(w7_61),.acc(r7_61),.res(r7_62),.clk(clk),.wout(w7_62));
	PE pe7_63(.x(x63),.w(w7_62),.acc(r7_62),.res(r7_63),.clk(clk),.wout(w7_63));
	PE pe7_64(.x(x64),.w(w7_63),.acc(r7_63),.res(r7_64),.clk(clk),.wout(w7_64));
	PE pe7_65(.x(x65),.w(w7_64),.acc(r7_64),.res(r7_65),.clk(clk),.wout(w7_65));
	PE pe7_66(.x(x66),.w(w7_65),.acc(r7_65),.res(r7_66),.clk(clk),.wout(w7_66));
	PE pe7_67(.x(x67),.w(w7_66),.acc(r7_66),.res(r7_67),.clk(clk),.wout(w7_67));
	PE pe7_68(.x(x68),.w(w7_67),.acc(r7_67),.res(r7_68),.clk(clk),.wout(w7_68));
	PE pe7_69(.x(x69),.w(w7_68),.acc(r7_68),.res(r7_69),.clk(clk),.wout(w7_69));
	PE pe7_70(.x(x70),.w(w7_69),.acc(r7_69),.res(r7_70),.clk(clk),.wout(w7_70));
	PE pe7_71(.x(x71),.w(w7_70),.acc(r7_70),.res(r7_71),.clk(clk),.wout(w7_71));
	PE pe7_72(.x(x72),.w(w7_71),.acc(r7_71),.res(r7_72),.clk(clk),.wout(w7_72));
	PE pe7_73(.x(x73),.w(w7_72),.acc(r7_72),.res(r7_73),.clk(clk),.wout(w7_73));
	PE pe7_74(.x(x74),.w(w7_73),.acc(r7_73),.res(r7_74),.clk(clk),.wout(w7_74));
	PE pe7_75(.x(x75),.w(w7_74),.acc(r7_74),.res(r7_75),.clk(clk),.wout(w7_75));
	PE pe7_76(.x(x76),.w(w7_75),.acc(r7_75),.res(r7_76),.clk(clk),.wout(w7_76));
	PE pe7_77(.x(x77),.w(w7_76),.acc(r7_76),.res(r7_77),.clk(clk),.wout(w7_77));
	PE pe7_78(.x(x78),.w(w7_77),.acc(r7_77),.res(r7_78),.clk(clk),.wout(w7_78));
	PE pe7_79(.x(x79),.w(w7_78),.acc(r7_78),.res(r7_79),.clk(clk),.wout(w7_79));
	PE pe7_80(.x(x80),.w(w7_79),.acc(r7_79),.res(r7_80),.clk(clk),.wout(w7_80));
	PE pe7_81(.x(x81),.w(w7_80),.acc(r7_80),.res(r7_81),.clk(clk),.wout(w7_81));
	PE pe7_82(.x(x82),.w(w7_81),.acc(r7_81),.res(r7_82),.clk(clk),.wout(w7_82));
	PE pe7_83(.x(x83),.w(w7_82),.acc(r7_82),.res(r7_83),.clk(clk),.wout(w7_83));
	PE pe7_84(.x(x84),.w(w7_83),.acc(r7_83),.res(r7_84),.clk(clk),.wout(w7_84));
	PE pe7_85(.x(x85),.w(w7_84),.acc(r7_84),.res(r7_85),.clk(clk),.wout(w7_85));
	PE pe7_86(.x(x86),.w(w7_85),.acc(r7_85),.res(r7_86),.clk(clk),.wout(w7_86));
	PE pe7_87(.x(x87),.w(w7_86),.acc(r7_86),.res(r7_87),.clk(clk),.wout(w7_87));
	PE pe7_88(.x(x88),.w(w7_87),.acc(r7_87),.res(r7_88),.clk(clk),.wout(w7_88));
	PE pe7_89(.x(x89),.w(w7_88),.acc(r7_88),.res(r7_89),.clk(clk),.wout(w7_89));
	PE pe7_90(.x(x90),.w(w7_89),.acc(r7_89),.res(r7_90),.clk(clk),.wout(w7_90));
	PE pe7_91(.x(x91),.w(w7_90),.acc(r7_90),.res(r7_91),.clk(clk),.wout(w7_91));
	PE pe7_92(.x(x92),.w(w7_91),.acc(r7_91),.res(r7_92),.clk(clk),.wout(w7_92));
	PE pe7_93(.x(x93),.w(w7_92),.acc(r7_92),.res(r7_93),.clk(clk),.wout(w7_93));
	PE pe7_94(.x(x94),.w(w7_93),.acc(r7_93),.res(r7_94),.clk(clk),.wout(w7_94));
	PE pe7_95(.x(x95),.w(w7_94),.acc(r7_94),.res(r7_95),.clk(clk),.wout(w7_95));
	PE pe7_96(.x(x96),.w(w7_95),.acc(r7_95),.res(r7_96),.clk(clk),.wout(w7_96));
	PE pe7_97(.x(x97),.w(w7_96),.acc(r7_96),.res(r7_97),.clk(clk),.wout(w7_97));
	PE pe7_98(.x(x98),.w(w7_97),.acc(r7_97),.res(r7_98),.clk(clk),.wout(w7_98));
	PE pe7_99(.x(x99),.w(w7_98),.acc(r7_98),.res(r7_99),.clk(clk),.wout(w7_99));
	PE pe7_100(.x(x100),.w(w7_99),.acc(r7_99),.res(r7_100),.clk(clk),.wout(w7_100));
	PE pe7_101(.x(x101),.w(w7_100),.acc(r7_100),.res(r7_101),.clk(clk),.wout(w7_101));
	PE pe7_102(.x(x102),.w(w7_101),.acc(r7_101),.res(r7_102),.clk(clk),.wout(w7_102));
	PE pe7_103(.x(x103),.w(w7_102),.acc(r7_102),.res(r7_103),.clk(clk),.wout(w7_103));
	PE pe7_104(.x(x104),.w(w7_103),.acc(r7_103),.res(r7_104),.clk(clk),.wout(w7_104));
	PE pe7_105(.x(x105),.w(w7_104),.acc(r7_104),.res(r7_105),.clk(clk),.wout(w7_105));
	PE pe7_106(.x(x106),.w(w7_105),.acc(r7_105),.res(r7_106),.clk(clk),.wout(w7_106));
	PE pe7_107(.x(x107),.w(w7_106),.acc(r7_106),.res(r7_107),.clk(clk),.wout(w7_107));
	PE pe7_108(.x(x108),.w(w7_107),.acc(r7_107),.res(r7_108),.clk(clk),.wout(w7_108));
	PE pe7_109(.x(x109),.w(w7_108),.acc(r7_108),.res(r7_109),.clk(clk),.wout(w7_109));
	PE pe7_110(.x(x110),.w(w7_109),.acc(r7_109),.res(r7_110),.clk(clk),.wout(w7_110));
	PE pe7_111(.x(x111),.w(w7_110),.acc(r7_110),.res(r7_111),.clk(clk),.wout(w7_111));
	PE pe7_112(.x(x112),.w(w7_111),.acc(r7_111),.res(r7_112),.clk(clk),.wout(w7_112));
	PE pe7_113(.x(x113),.w(w7_112),.acc(r7_112),.res(r7_113),.clk(clk),.wout(w7_113));
	PE pe7_114(.x(x114),.w(w7_113),.acc(r7_113),.res(r7_114),.clk(clk),.wout(w7_114));
	PE pe7_115(.x(x115),.w(w7_114),.acc(r7_114),.res(r7_115),.clk(clk),.wout(w7_115));
	PE pe7_116(.x(x116),.w(w7_115),.acc(r7_115),.res(r7_116),.clk(clk),.wout(w7_116));
	PE pe7_117(.x(x117),.w(w7_116),.acc(r7_116),.res(r7_117),.clk(clk),.wout(w7_117));
	PE pe7_118(.x(x118),.w(w7_117),.acc(r7_117),.res(r7_118),.clk(clk),.wout(w7_118));
	PE pe7_119(.x(x119),.w(w7_118),.acc(r7_118),.res(r7_119),.clk(clk),.wout(w7_119));
	PE pe7_120(.x(x120),.w(w7_119),.acc(r7_119),.res(r7_120),.clk(clk),.wout(w7_120));
	PE pe7_121(.x(x121),.w(w7_120),.acc(r7_120),.res(r7_121),.clk(clk),.wout(w7_121));
	PE pe7_122(.x(x122),.w(w7_121),.acc(r7_121),.res(r7_122),.clk(clk),.wout(w7_122));
	PE pe7_123(.x(x123),.w(w7_122),.acc(r7_122),.res(r7_123),.clk(clk),.wout(w7_123));
	PE pe7_124(.x(x124),.w(w7_123),.acc(r7_123),.res(r7_124),.clk(clk),.wout(w7_124));
	PE pe7_125(.x(x125),.w(w7_124),.acc(r7_124),.res(r7_125),.clk(clk),.wout(w7_125));
	PE pe7_126(.x(x126),.w(w7_125),.acc(r7_125),.res(r7_126),.clk(clk),.wout(w7_126));
	PE pe7_127(.x(x127),.w(w7_126),.acc(r7_126),.res(result7),.clk(clk),.wout(weight7));

	PE pe8_0(.x(x0),.w(w8),.acc(32'h0),.res(r8_0),.clk(clk),.wout(w8_0));
	PE pe8_1(.x(x1),.w(w8_0),.acc(r8_0),.res(r8_1),.clk(clk),.wout(w8_1));
	PE pe8_2(.x(x2),.w(w8_1),.acc(r8_1),.res(r8_2),.clk(clk),.wout(w8_2));
	PE pe8_3(.x(x3),.w(w8_2),.acc(r8_2),.res(r8_3),.clk(clk),.wout(w8_3));
	PE pe8_4(.x(x4),.w(w8_3),.acc(r8_3),.res(r8_4),.clk(clk),.wout(w8_4));
	PE pe8_5(.x(x5),.w(w8_4),.acc(r8_4),.res(r8_5),.clk(clk),.wout(w8_5));
	PE pe8_6(.x(x6),.w(w8_5),.acc(r8_5),.res(r8_6),.clk(clk),.wout(w8_6));
	PE pe8_7(.x(x7),.w(w8_6),.acc(r8_6),.res(r8_7),.clk(clk),.wout(w8_7));
	PE pe8_8(.x(x8),.w(w8_7),.acc(r8_7),.res(r8_8),.clk(clk),.wout(w8_8));
	PE pe8_9(.x(x9),.w(w8_8),.acc(r8_8),.res(r8_9),.clk(clk),.wout(w8_9));
	PE pe8_10(.x(x10),.w(w8_9),.acc(r8_9),.res(r8_10),.clk(clk),.wout(w8_10));
	PE pe8_11(.x(x11),.w(w8_10),.acc(r8_10),.res(r8_11),.clk(clk),.wout(w8_11));
	PE pe8_12(.x(x12),.w(w8_11),.acc(r8_11),.res(r8_12),.clk(clk),.wout(w8_12));
	PE pe8_13(.x(x13),.w(w8_12),.acc(r8_12),.res(r8_13),.clk(clk),.wout(w8_13));
	PE pe8_14(.x(x14),.w(w8_13),.acc(r8_13),.res(r8_14),.clk(clk),.wout(w8_14));
	PE pe8_15(.x(x15),.w(w8_14),.acc(r8_14),.res(r8_15),.clk(clk),.wout(w8_15));
	PE pe8_16(.x(x16),.w(w8_15),.acc(r8_15),.res(r8_16),.clk(clk),.wout(w8_16));
	PE pe8_17(.x(x17),.w(w8_16),.acc(r8_16),.res(r8_17),.clk(clk),.wout(w8_17));
	PE pe8_18(.x(x18),.w(w8_17),.acc(r8_17),.res(r8_18),.clk(clk),.wout(w8_18));
	PE pe8_19(.x(x19),.w(w8_18),.acc(r8_18),.res(r8_19),.clk(clk),.wout(w8_19));
	PE pe8_20(.x(x20),.w(w8_19),.acc(r8_19),.res(r8_20),.clk(clk),.wout(w8_20));
	PE pe8_21(.x(x21),.w(w8_20),.acc(r8_20),.res(r8_21),.clk(clk),.wout(w8_21));
	PE pe8_22(.x(x22),.w(w8_21),.acc(r8_21),.res(r8_22),.clk(clk),.wout(w8_22));
	PE pe8_23(.x(x23),.w(w8_22),.acc(r8_22),.res(r8_23),.clk(clk),.wout(w8_23));
	PE pe8_24(.x(x24),.w(w8_23),.acc(r8_23),.res(r8_24),.clk(clk),.wout(w8_24));
	PE pe8_25(.x(x25),.w(w8_24),.acc(r8_24),.res(r8_25),.clk(clk),.wout(w8_25));
	PE pe8_26(.x(x26),.w(w8_25),.acc(r8_25),.res(r8_26),.clk(clk),.wout(w8_26));
	PE pe8_27(.x(x27),.w(w8_26),.acc(r8_26),.res(r8_27),.clk(clk),.wout(w8_27));
	PE pe8_28(.x(x28),.w(w8_27),.acc(r8_27),.res(r8_28),.clk(clk),.wout(w8_28));
	PE pe8_29(.x(x29),.w(w8_28),.acc(r8_28),.res(r8_29),.clk(clk),.wout(w8_29));
	PE pe8_30(.x(x30),.w(w8_29),.acc(r8_29),.res(r8_30),.clk(clk),.wout(w8_30));
	PE pe8_31(.x(x31),.w(w8_30),.acc(r8_30),.res(r8_31),.clk(clk),.wout(w8_31));
	PE pe8_32(.x(x32),.w(w8_31),.acc(r8_31),.res(r8_32),.clk(clk),.wout(w8_32));
	PE pe8_33(.x(x33),.w(w8_32),.acc(r8_32),.res(r8_33),.clk(clk),.wout(w8_33));
	PE pe8_34(.x(x34),.w(w8_33),.acc(r8_33),.res(r8_34),.clk(clk),.wout(w8_34));
	PE pe8_35(.x(x35),.w(w8_34),.acc(r8_34),.res(r8_35),.clk(clk),.wout(w8_35));
	PE pe8_36(.x(x36),.w(w8_35),.acc(r8_35),.res(r8_36),.clk(clk),.wout(w8_36));
	PE pe8_37(.x(x37),.w(w8_36),.acc(r8_36),.res(r8_37),.clk(clk),.wout(w8_37));
	PE pe8_38(.x(x38),.w(w8_37),.acc(r8_37),.res(r8_38),.clk(clk),.wout(w8_38));
	PE pe8_39(.x(x39),.w(w8_38),.acc(r8_38),.res(r8_39),.clk(clk),.wout(w8_39));
	PE pe8_40(.x(x40),.w(w8_39),.acc(r8_39),.res(r8_40),.clk(clk),.wout(w8_40));
	PE pe8_41(.x(x41),.w(w8_40),.acc(r8_40),.res(r8_41),.clk(clk),.wout(w8_41));
	PE pe8_42(.x(x42),.w(w8_41),.acc(r8_41),.res(r8_42),.clk(clk),.wout(w8_42));
	PE pe8_43(.x(x43),.w(w8_42),.acc(r8_42),.res(r8_43),.clk(clk),.wout(w8_43));
	PE pe8_44(.x(x44),.w(w8_43),.acc(r8_43),.res(r8_44),.clk(clk),.wout(w8_44));
	PE pe8_45(.x(x45),.w(w8_44),.acc(r8_44),.res(r8_45),.clk(clk),.wout(w8_45));
	PE pe8_46(.x(x46),.w(w8_45),.acc(r8_45),.res(r8_46),.clk(clk),.wout(w8_46));
	PE pe8_47(.x(x47),.w(w8_46),.acc(r8_46),.res(r8_47),.clk(clk),.wout(w8_47));
	PE pe8_48(.x(x48),.w(w8_47),.acc(r8_47),.res(r8_48),.clk(clk),.wout(w8_48));
	PE pe8_49(.x(x49),.w(w8_48),.acc(r8_48),.res(r8_49),.clk(clk),.wout(w8_49));
	PE pe8_50(.x(x50),.w(w8_49),.acc(r8_49),.res(r8_50),.clk(clk),.wout(w8_50));
	PE pe8_51(.x(x51),.w(w8_50),.acc(r8_50),.res(r8_51),.clk(clk),.wout(w8_51));
	PE pe8_52(.x(x52),.w(w8_51),.acc(r8_51),.res(r8_52),.clk(clk),.wout(w8_52));
	PE pe8_53(.x(x53),.w(w8_52),.acc(r8_52),.res(r8_53),.clk(clk),.wout(w8_53));
	PE pe8_54(.x(x54),.w(w8_53),.acc(r8_53),.res(r8_54),.clk(clk),.wout(w8_54));
	PE pe8_55(.x(x55),.w(w8_54),.acc(r8_54),.res(r8_55),.clk(clk),.wout(w8_55));
	PE pe8_56(.x(x56),.w(w8_55),.acc(r8_55),.res(r8_56),.clk(clk),.wout(w8_56));
	PE pe8_57(.x(x57),.w(w8_56),.acc(r8_56),.res(r8_57),.clk(clk),.wout(w8_57));
	PE pe8_58(.x(x58),.w(w8_57),.acc(r8_57),.res(r8_58),.clk(clk),.wout(w8_58));
	PE pe8_59(.x(x59),.w(w8_58),.acc(r8_58),.res(r8_59),.clk(clk),.wout(w8_59));
	PE pe8_60(.x(x60),.w(w8_59),.acc(r8_59),.res(r8_60),.clk(clk),.wout(w8_60));
	PE pe8_61(.x(x61),.w(w8_60),.acc(r8_60),.res(r8_61),.clk(clk),.wout(w8_61));
	PE pe8_62(.x(x62),.w(w8_61),.acc(r8_61),.res(r8_62),.clk(clk),.wout(w8_62));
	PE pe8_63(.x(x63),.w(w8_62),.acc(r8_62),.res(r8_63),.clk(clk),.wout(w8_63));
	PE pe8_64(.x(x64),.w(w8_63),.acc(r8_63),.res(r8_64),.clk(clk),.wout(w8_64));
	PE pe8_65(.x(x65),.w(w8_64),.acc(r8_64),.res(r8_65),.clk(clk),.wout(w8_65));
	PE pe8_66(.x(x66),.w(w8_65),.acc(r8_65),.res(r8_66),.clk(clk),.wout(w8_66));
	PE pe8_67(.x(x67),.w(w8_66),.acc(r8_66),.res(r8_67),.clk(clk),.wout(w8_67));
	PE pe8_68(.x(x68),.w(w8_67),.acc(r8_67),.res(r8_68),.clk(clk),.wout(w8_68));
	PE pe8_69(.x(x69),.w(w8_68),.acc(r8_68),.res(r8_69),.clk(clk),.wout(w8_69));
	PE pe8_70(.x(x70),.w(w8_69),.acc(r8_69),.res(r8_70),.clk(clk),.wout(w8_70));
	PE pe8_71(.x(x71),.w(w8_70),.acc(r8_70),.res(r8_71),.clk(clk),.wout(w8_71));
	PE pe8_72(.x(x72),.w(w8_71),.acc(r8_71),.res(r8_72),.clk(clk),.wout(w8_72));
	PE pe8_73(.x(x73),.w(w8_72),.acc(r8_72),.res(r8_73),.clk(clk),.wout(w8_73));
	PE pe8_74(.x(x74),.w(w8_73),.acc(r8_73),.res(r8_74),.clk(clk),.wout(w8_74));
	PE pe8_75(.x(x75),.w(w8_74),.acc(r8_74),.res(r8_75),.clk(clk),.wout(w8_75));
	PE pe8_76(.x(x76),.w(w8_75),.acc(r8_75),.res(r8_76),.clk(clk),.wout(w8_76));
	PE pe8_77(.x(x77),.w(w8_76),.acc(r8_76),.res(r8_77),.clk(clk),.wout(w8_77));
	PE pe8_78(.x(x78),.w(w8_77),.acc(r8_77),.res(r8_78),.clk(clk),.wout(w8_78));
	PE pe8_79(.x(x79),.w(w8_78),.acc(r8_78),.res(r8_79),.clk(clk),.wout(w8_79));
	PE pe8_80(.x(x80),.w(w8_79),.acc(r8_79),.res(r8_80),.clk(clk),.wout(w8_80));
	PE pe8_81(.x(x81),.w(w8_80),.acc(r8_80),.res(r8_81),.clk(clk),.wout(w8_81));
	PE pe8_82(.x(x82),.w(w8_81),.acc(r8_81),.res(r8_82),.clk(clk),.wout(w8_82));
	PE pe8_83(.x(x83),.w(w8_82),.acc(r8_82),.res(r8_83),.clk(clk),.wout(w8_83));
	PE pe8_84(.x(x84),.w(w8_83),.acc(r8_83),.res(r8_84),.clk(clk),.wout(w8_84));
	PE pe8_85(.x(x85),.w(w8_84),.acc(r8_84),.res(r8_85),.clk(clk),.wout(w8_85));
	PE pe8_86(.x(x86),.w(w8_85),.acc(r8_85),.res(r8_86),.clk(clk),.wout(w8_86));
	PE pe8_87(.x(x87),.w(w8_86),.acc(r8_86),.res(r8_87),.clk(clk),.wout(w8_87));
	PE pe8_88(.x(x88),.w(w8_87),.acc(r8_87),.res(r8_88),.clk(clk),.wout(w8_88));
	PE pe8_89(.x(x89),.w(w8_88),.acc(r8_88),.res(r8_89),.clk(clk),.wout(w8_89));
	PE pe8_90(.x(x90),.w(w8_89),.acc(r8_89),.res(r8_90),.clk(clk),.wout(w8_90));
	PE pe8_91(.x(x91),.w(w8_90),.acc(r8_90),.res(r8_91),.clk(clk),.wout(w8_91));
	PE pe8_92(.x(x92),.w(w8_91),.acc(r8_91),.res(r8_92),.clk(clk),.wout(w8_92));
	PE pe8_93(.x(x93),.w(w8_92),.acc(r8_92),.res(r8_93),.clk(clk),.wout(w8_93));
	PE pe8_94(.x(x94),.w(w8_93),.acc(r8_93),.res(r8_94),.clk(clk),.wout(w8_94));
	PE pe8_95(.x(x95),.w(w8_94),.acc(r8_94),.res(r8_95),.clk(clk),.wout(w8_95));
	PE pe8_96(.x(x96),.w(w8_95),.acc(r8_95),.res(r8_96),.clk(clk),.wout(w8_96));
	PE pe8_97(.x(x97),.w(w8_96),.acc(r8_96),.res(r8_97),.clk(clk),.wout(w8_97));
	PE pe8_98(.x(x98),.w(w8_97),.acc(r8_97),.res(r8_98),.clk(clk),.wout(w8_98));
	PE pe8_99(.x(x99),.w(w8_98),.acc(r8_98),.res(r8_99),.clk(clk),.wout(w8_99));
	PE pe8_100(.x(x100),.w(w8_99),.acc(r8_99),.res(r8_100),.clk(clk),.wout(w8_100));
	PE pe8_101(.x(x101),.w(w8_100),.acc(r8_100),.res(r8_101),.clk(clk),.wout(w8_101));
	PE pe8_102(.x(x102),.w(w8_101),.acc(r8_101),.res(r8_102),.clk(clk),.wout(w8_102));
	PE pe8_103(.x(x103),.w(w8_102),.acc(r8_102),.res(r8_103),.clk(clk),.wout(w8_103));
	PE pe8_104(.x(x104),.w(w8_103),.acc(r8_103),.res(r8_104),.clk(clk),.wout(w8_104));
	PE pe8_105(.x(x105),.w(w8_104),.acc(r8_104),.res(r8_105),.clk(clk),.wout(w8_105));
	PE pe8_106(.x(x106),.w(w8_105),.acc(r8_105),.res(r8_106),.clk(clk),.wout(w8_106));
	PE pe8_107(.x(x107),.w(w8_106),.acc(r8_106),.res(r8_107),.clk(clk),.wout(w8_107));
	PE pe8_108(.x(x108),.w(w8_107),.acc(r8_107),.res(r8_108),.clk(clk),.wout(w8_108));
	PE pe8_109(.x(x109),.w(w8_108),.acc(r8_108),.res(r8_109),.clk(clk),.wout(w8_109));
	PE pe8_110(.x(x110),.w(w8_109),.acc(r8_109),.res(r8_110),.clk(clk),.wout(w8_110));
	PE pe8_111(.x(x111),.w(w8_110),.acc(r8_110),.res(r8_111),.clk(clk),.wout(w8_111));
	PE pe8_112(.x(x112),.w(w8_111),.acc(r8_111),.res(r8_112),.clk(clk),.wout(w8_112));
	PE pe8_113(.x(x113),.w(w8_112),.acc(r8_112),.res(r8_113),.clk(clk),.wout(w8_113));
	PE pe8_114(.x(x114),.w(w8_113),.acc(r8_113),.res(r8_114),.clk(clk),.wout(w8_114));
	PE pe8_115(.x(x115),.w(w8_114),.acc(r8_114),.res(r8_115),.clk(clk),.wout(w8_115));
	PE pe8_116(.x(x116),.w(w8_115),.acc(r8_115),.res(r8_116),.clk(clk),.wout(w8_116));
	PE pe8_117(.x(x117),.w(w8_116),.acc(r8_116),.res(r8_117),.clk(clk),.wout(w8_117));
	PE pe8_118(.x(x118),.w(w8_117),.acc(r8_117),.res(r8_118),.clk(clk),.wout(w8_118));
	PE pe8_119(.x(x119),.w(w8_118),.acc(r8_118),.res(r8_119),.clk(clk),.wout(w8_119));
	PE pe8_120(.x(x120),.w(w8_119),.acc(r8_119),.res(r8_120),.clk(clk),.wout(w8_120));
	PE pe8_121(.x(x121),.w(w8_120),.acc(r8_120),.res(r8_121),.clk(clk),.wout(w8_121));
	PE pe8_122(.x(x122),.w(w8_121),.acc(r8_121),.res(r8_122),.clk(clk),.wout(w8_122));
	PE pe8_123(.x(x123),.w(w8_122),.acc(r8_122),.res(r8_123),.clk(clk),.wout(w8_123));
	PE pe8_124(.x(x124),.w(w8_123),.acc(r8_123),.res(r8_124),.clk(clk),.wout(w8_124));
	PE pe8_125(.x(x125),.w(w8_124),.acc(r8_124),.res(r8_125),.clk(clk),.wout(w8_125));
	PE pe8_126(.x(x126),.w(w8_125),.acc(r8_125),.res(r8_126),.clk(clk),.wout(w8_126));
	PE pe8_127(.x(x127),.w(w8_126),.acc(r8_126),.res(result8),.clk(clk),.wout(weight8));

	PE pe9_0(.x(x0),.w(w9),.acc(32'h0),.res(r9_0),.clk(clk),.wout(w9_0));
	PE pe9_1(.x(x1),.w(w9_0),.acc(r9_0),.res(r9_1),.clk(clk),.wout(w9_1));
	PE pe9_2(.x(x2),.w(w9_1),.acc(r9_1),.res(r9_2),.clk(clk),.wout(w9_2));
	PE pe9_3(.x(x3),.w(w9_2),.acc(r9_2),.res(r9_3),.clk(clk),.wout(w9_3));
	PE pe9_4(.x(x4),.w(w9_3),.acc(r9_3),.res(r9_4),.clk(clk),.wout(w9_4));
	PE pe9_5(.x(x5),.w(w9_4),.acc(r9_4),.res(r9_5),.clk(clk),.wout(w9_5));
	PE pe9_6(.x(x6),.w(w9_5),.acc(r9_5),.res(r9_6),.clk(clk),.wout(w9_6));
	PE pe9_7(.x(x7),.w(w9_6),.acc(r9_6),.res(r9_7),.clk(clk),.wout(w9_7));
	PE pe9_8(.x(x8),.w(w9_7),.acc(r9_7),.res(r9_8),.clk(clk),.wout(w9_8));
	PE pe9_9(.x(x9),.w(w9_8),.acc(r9_8),.res(r9_9),.clk(clk),.wout(w9_9));
	PE pe9_10(.x(x10),.w(w9_9),.acc(r9_9),.res(r9_10),.clk(clk),.wout(w9_10));
	PE pe9_11(.x(x11),.w(w9_10),.acc(r9_10),.res(r9_11),.clk(clk),.wout(w9_11));
	PE pe9_12(.x(x12),.w(w9_11),.acc(r9_11),.res(r9_12),.clk(clk),.wout(w9_12));
	PE pe9_13(.x(x13),.w(w9_12),.acc(r9_12),.res(r9_13),.clk(clk),.wout(w9_13));
	PE pe9_14(.x(x14),.w(w9_13),.acc(r9_13),.res(r9_14),.clk(clk),.wout(w9_14));
	PE pe9_15(.x(x15),.w(w9_14),.acc(r9_14),.res(r9_15),.clk(clk),.wout(w9_15));
	PE pe9_16(.x(x16),.w(w9_15),.acc(r9_15),.res(r9_16),.clk(clk),.wout(w9_16));
	PE pe9_17(.x(x17),.w(w9_16),.acc(r9_16),.res(r9_17),.clk(clk),.wout(w9_17));
	PE pe9_18(.x(x18),.w(w9_17),.acc(r9_17),.res(r9_18),.clk(clk),.wout(w9_18));
	PE pe9_19(.x(x19),.w(w9_18),.acc(r9_18),.res(r9_19),.clk(clk),.wout(w9_19));
	PE pe9_20(.x(x20),.w(w9_19),.acc(r9_19),.res(r9_20),.clk(clk),.wout(w9_20));
	PE pe9_21(.x(x21),.w(w9_20),.acc(r9_20),.res(r9_21),.clk(clk),.wout(w9_21));
	PE pe9_22(.x(x22),.w(w9_21),.acc(r9_21),.res(r9_22),.clk(clk),.wout(w9_22));
	PE pe9_23(.x(x23),.w(w9_22),.acc(r9_22),.res(r9_23),.clk(clk),.wout(w9_23));
	PE pe9_24(.x(x24),.w(w9_23),.acc(r9_23),.res(r9_24),.clk(clk),.wout(w9_24));
	PE pe9_25(.x(x25),.w(w9_24),.acc(r9_24),.res(r9_25),.clk(clk),.wout(w9_25));
	PE pe9_26(.x(x26),.w(w9_25),.acc(r9_25),.res(r9_26),.clk(clk),.wout(w9_26));
	PE pe9_27(.x(x27),.w(w9_26),.acc(r9_26),.res(r9_27),.clk(clk),.wout(w9_27));
	PE pe9_28(.x(x28),.w(w9_27),.acc(r9_27),.res(r9_28),.clk(clk),.wout(w9_28));
	PE pe9_29(.x(x29),.w(w9_28),.acc(r9_28),.res(r9_29),.clk(clk),.wout(w9_29));
	PE pe9_30(.x(x30),.w(w9_29),.acc(r9_29),.res(r9_30),.clk(clk),.wout(w9_30));
	PE pe9_31(.x(x31),.w(w9_30),.acc(r9_30),.res(r9_31),.clk(clk),.wout(w9_31));
	PE pe9_32(.x(x32),.w(w9_31),.acc(r9_31),.res(r9_32),.clk(clk),.wout(w9_32));
	PE pe9_33(.x(x33),.w(w9_32),.acc(r9_32),.res(r9_33),.clk(clk),.wout(w9_33));
	PE pe9_34(.x(x34),.w(w9_33),.acc(r9_33),.res(r9_34),.clk(clk),.wout(w9_34));
	PE pe9_35(.x(x35),.w(w9_34),.acc(r9_34),.res(r9_35),.clk(clk),.wout(w9_35));
	PE pe9_36(.x(x36),.w(w9_35),.acc(r9_35),.res(r9_36),.clk(clk),.wout(w9_36));
	PE pe9_37(.x(x37),.w(w9_36),.acc(r9_36),.res(r9_37),.clk(clk),.wout(w9_37));
	PE pe9_38(.x(x38),.w(w9_37),.acc(r9_37),.res(r9_38),.clk(clk),.wout(w9_38));
	PE pe9_39(.x(x39),.w(w9_38),.acc(r9_38),.res(r9_39),.clk(clk),.wout(w9_39));
	PE pe9_40(.x(x40),.w(w9_39),.acc(r9_39),.res(r9_40),.clk(clk),.wout(w9_40));
	PE pe9_41(.x(x41),.w(w9_40),.acc(r9_40),.res(r9_41),.clk(clk),.wout(w9_41));
	PE pe9_42(.x(x42),.w(w9_41),.acc(r9_41),.res(r9_42),.clk(clk),.wout(w9_42));
	PE pe9_43(.x(x43),.w(w9_42),.acc(r9_42),.res(r9_43),.clk(clk),.wout(w9_43));
	PE pe9_44(.x(x44),.w(w9_43),.acc(r9_43),.res(r9_44),.clk(clk),.wout(w9_44));
	PE pe9_45(.x(x45),.w(w9_44),.acc(r9_44),.res(r9_45),.clk(clk),.wout(w9_45));
	PE pe9_46(.x(x46),.w(w9_45),.acc(r9_45),.res(r9_46),.clk(clk),.wout(w9_46));
	PE pe9_47(.x(x47),.w(w9_46),.acc(r9_46),.res(r9_47),.clk(clk),.wout(w9_47));
	PE pe9_48(.x(x48),.w(w9_47),.acc(r9_47),.res(r9_48),.clk(clk),.wout(w9_48));
	PE pe9_49(.x(x49),.w(w9_48),.acc(r9_48),.res(r9_49),.clk(clk),.wout(w9_49));
	PE pe9_50(.x(x50),.w(w9_49),.acc(r9_49),.res(r9_50),.clk(clk),.wout(w9_50));
	PE pe9_51(.x(x51),.w(w9_50),.acc(r9_50),.res(r9_51),.clk(clk),.wout(w9_51));
	PE pe9_52(.x(x52),.w(w9_51),.acc(r9_51),.res(r9_52),.clk(clk),.wout(w9_52));
	PE pe9_53(.x(x53),.w(w9_52),.acc(r9_52),.res(r9_53),.clk(clk),.wout(w9_53));
	PE pe9_54(.x(x54),.w(w9_53),.acc(r9_53),.res(r9_54),.clk(clk),.wout(w9_54));
	PE pe9_55(.x(x55),.w(w9_54),.acc(r9_54),.res(r9_55),.clk(clk),.wout(w9_55));
	PE pe9_56(.x(x56),.w(w9_55),.acc(r9_55),.res(r9_56),.clk(clk),.wout(w9_56));
	PE pe9_57(.x(x57),.w(w9_56),.acc(r9_56),.res(r9_57),.clk(clk),.wout(w9_57));
	PE pe9_58(.x(x58),.w(w9_57),.acc(r9_57),.res(r9_58),.clk(clk),.wout(w9_58));
	PE pe9_59(.x(x59),.w(w9_58),.acc(r9_58),.res(r9_59),.clk(clk),.wout(w9_59));
	PE pe9_60(.x(x60),.w(w9_59),.acc(r9_59),.res(r9_60),.clk(clk),.wout(w9_60));
	PE pe9_61(.x(x61),.w(w9_60),.acc(r9_60),.res(r9_61),.clk(clk),.wout(w9_61));
	PE pe9_62(.x(x62),.w(w9_61),.acc(r9_61),.res(r9_62),.clk(clk),.wout(w9_62));
	PE pe9_63(.x(x63),.w(w9_62),.acc(r9_62),.res(r9_63),.clk(clk),.wout(w9_63));
	PE pe9_64(.x(x64),.w(w9_63),.acc(r9_63),.res(r9_64),.clk(clk),.wout(w9_64));
	PE pe9_65(.x(x65),.w(w9_64),.acc(r9_64),.res(r9_65),.clk(clk),.wout(w9_65));
	PE pe9_66(.x(x66),.w(w9_65),.acc(r9_65),.res(r9_66),.clk(clk),.wout(w9_66));
	PE pe9_67(.x(x67),.w(w9_66),.acc(r9_66),.res(r9_67),.clk(clk),.wout(w9_67));
	PE pe9_68(.x(x68),.w(w9_67),.acc(r9_67),.res(r9_68),.clk(clk),.wout(w9_68));
	PE pe9_69(.x(x69),.w(w9_68),.acc(r9_68),.res(r9_69),.clk(clk),.wout(w9_69));
	PE pe9_70(.x(x70),.w(w9_69),.acc(r9_69),.res(r9_70),.clk(clk),.wout(w9_70));
	PE pe9_71(.x(x71),.w(w9_70),.acc(r9_70),.res(r9_71),.clk(clk),.wout(w9_71));
	PE pe9_72(.x(x72),.w(w9_71),.acc(r9_71),.res(r9_72),.clk(clk),.wout(w9_72));
	PE pe9_73(.x(x73),.w(w9_72),.acc(r9_72),.res(r9_73),.clk(clk),.wout(w9_73));
	PE pe9_74(.x(x74),.w(w9_73),.acc(r9_73),.res(r9_74),.clk(clk),.wout(w9_74));
	PE pe9_75(.x(x75),.w(w9_74),.acc(r9_74),.res(r9_75),.clk(clk),.wout(w9_75));
	PE pe9_76(.x(x76),.w(w9_75),.acc(r9_75),.res(r9_76),.clk(clk),.wout(w9_76));
	PE pe9_77(.x(x77),.w(w9_76),.acc(r9_76),.res(r9_77),.clk(clk),.wout(w9_77));
	PE pe9_78(.x(x78),.w(w9_77),.acc(r9_77),.res(r9_78),.clk(clk),.wout(w9_78));
	PE pe9_79(.x(x79),.w(w9_78),.acc(r9_78),.res(r9_79),.clk(clk),.wout(w9_79));
	PE pe9_80(.x(x80),.w(w9_79),.acc(r9_79),.res(r9_80),.clk(clk),.wout(w9_80));
	PE pe9_81(.x(x81),.w(w9_80),.acc(r9_80),.res(r9_81),.clk(clk),.wout(w9_81));
	PE pe9_82(.x(x82),.w(w9_81),.acc(r9_81),.res(r9_82),.clk(clk),.wout(w9_82));
	PE pe9_83(.x(x83),.w(w9_82),.acc(r9_82),.res(r9_83),.clk(clk),.wout(w9_83));
	PE pe9_84(.x(x84),.w(w9_83),.acc(r9_83),.res(r9_84),.clk(clk),.wout(w9_84));
	PE pe9_85(.x(x85),.w(w9_84),.acc(r9_84),.res(r9_85),.clk(clk),.wout(w9_85));
	PE pe9_86(.x(x86),.w(w9_85),.acc(r9_85),.res(r9_86),.clk(clk),.wout(w9_86));
	PE pe9_87(.x(x87),.w(w9_86),.acc(r9_86),.res(r9_87),.clk(clk),.wout(w9_87));
	PE pe9_88(.x(x88),.w(w9_87),.acc(r9_87),.res(r9_88),.clk(clk),.wout(w9_88));
	PE pe9_89(.x(x89),.w(w9_88),.acc(r9_88),.res(r9_89),.clk(clk),.wout(w9_89));
	PE pe9_90(.x(x90),.w(w9_89),.acc(r9_89),.res(r9_90),.clk(clk),.wout(w9_90));
	PE pe9_91(.x(x91),.w(w9_90),.acc(r9_90),.res(r9_91),.clk(clk),.wout(w9_91));
	PE pe9_92(.x(x92),.w(w9_91),.acc(r9_91),.res(r9_92),.clk(clk),.wout(w9_92));
	PE pe9_93(.x(x93),.w(w9_92),.acc(r9_92),.res(r9_93),.clk(clk),.wout(w9_93));
	PE pe9_94(.x(x94),.w(w9_93),.acc(r9_93),.res(r9_94),.clk(clk),.wout(w9_94));
	PE pe9_95(.x(x95),.w(w9_94),.acc(r9_94),.res(r9_95),.clk(clk),.wout(w9_95));
	PE pe9_96(.x(x96),.w(w9_95),.acc(r9_95),.res(r9_96),.clk(clk),.wout(w9_96));
	PE pe9_97(.x(x97),.w(w9_96),.acc(r9_96),.res(r9_97),.clk(clk),.wout(w9_97));
	PE pe9_98(.x(x98),.w(w9_97),.acc(r9_97),.res(r9_98),.clk(clk),.wout(w9_98));
	PE pe9_99(.x(x99),.w(w9_98),.acc(r9_98),.res(r9_99),.clk(clk),.wout(w9_99));
	PE pe9_100(.x(x100),.w(w9_99),.acc(r9_99),.res(r9_100),.clk(clk),.wout(w9_100));
	PE pe9_101(.x(x101),.w(w9_100),.acc(r9_100),.res(r9_101),.clk(clk),.wout(w9_101));
	PE pe9_102(.x(x102),.w(w9_101),.acc(r9_101),.res(r9_102),.clk(clk),.wout(w9_102));
	PE pe9_103(.x(x103),.w(w9_102),.acc(r9_102),.res(r9_103),.clk(clk),.wout(w9_103));
	PE pe9_104(.x(x104),.w(w9_103),.acc(r9_103),.res(r9_104),.clk(clk),.wout(w9_104));
	PE pe9_105(.x(x105),.w(w9_104),.acc(r9_104),.res(r9_105),.clk(clk),.wout(w9_105));
	PE pe9_106(.x(x106),.w(w9_105),.acc(r9_105),.res(r9_106),.clk(clk),.wout(w9_106));
	PE pe9_107(.x(x107),.w(w9_106),.acc(r9_106),.res(r9_107),.clk(clk),.wout(w9_107));
	PE pe9_108(.x(x108),.w(w9_107),.acc(r9_107),.res(r9_108),.clk(clk),.wout(w9_108));
	PE pe9_109(.x(x109),.w(w9_108),.acc(r9_108),.res(r9_109),.clk(clk),.wout(w9_109));
	PE pe9_110(.x(x110),.w(w9_109),.acc(r9_109),.res(r9_110),.clk(clk),.wout(w9_110));
	PE pe9_111(.x(x111),.w(w9_110),.acc(r9_110),.res(r9_111),.clk(clk),.wout(w9_111));
	PE pe9_112(.x(x112),.w(w9_111),.acc(r9_111),.res(r9_112),.clk(clk),.wout(w9_112));
	PE pe9_113(.x(x113),.w(w9_112),.acc(r9_112),.res(r9_113),.clk(clk),.wout(w9_113));
	PE pe9_114(.x(x114),.w(w9_113),.acc(r9_113),.res(r9_114),.clk(clk),.wout(w9_114));
	PE pe9_115(.x(x115),.w(w9_114),.acc(r9_114),.res(r9_115),.clk(clk),.wout(w9_115));
	PE pe9_116(.x(x116),.w(w9_115),.acc(r9_115),.res(r9_116),.clk(clk),.wout(w9_116));
	PE pe9_117(.x(x117),.w(w9_116),.acc(r9_116),.res(r9_117),.clk(clk),.wout(w9_117));
	PE pe9_118(.x(x118),.w(w9_117),.acc(r9_117),.res(r9_118),.clk(clk),.wout(w9_118));
	PE pe9_119(.x(x119),.w(w9_118),.acc(r9_118),.res(r9_119),.clk(clk),.wout(w9_119));
	PE pe9_120(.x(x120),.w(w9_119),.acc(r9_119),.res(r9_120),.clk(clk),.wout(w9_120));
	PE pe9_121(.x(x121),.w(w9_120),.acc(r9_120),.res(r9_121),.clk(clk),.wout(w9_121));
	PE pe9_122(.x(x122),.w(w9_121),.acc(r9_121),.res(r9_122),.clk(clk),.wout(w9_122));
	PE pe9_123(.x(x123),.w(w9_122),.acc(r9_122),.res(r9_123),.clk(clk),.wout(w9_123));
	PE pe9_124(.x(x124),.w(w9_123),.acc(r9_123),.res(r9_124),.clk(clk),.wout(w9_124));
	PE pe9_125(.x(x125),.w(w9_124),.acc(r9_124),.res(r9_125),.clk(clk),.wout(w9_125));
	PE pe9_126(.x(x126),.w(w9_125),.acc(r9_125),.res(r9_126),.clk(clk),.wout(w9_126));
	PE pe9_127(.x(x127),.w(w9_126),.acc(r9_126),.res(result9),.clk(clk),.wout(weight9));

	PE pe10_0(.x(x0),.w(w10),.acc(32'h0),.res(r10_0),.clk(clk),.wout(w10_0));
	PE pe10_1(.x(x1),.w(w10_0),.acc(r10_0),.res(r10_1),.clk(clk),.wout(w10_1));
	PE pe10_2(.x(x2),.w(w10_1),.acc(r10_1),.res(r10_2),.clk(clk),.wout(w10_2));
	PE pe10_3(.x(x3),.w(w10_2),.acc(r10_2),.res(r10_3),.clk(clk),.wout(w10_3));
	PE pe10_4(.x(x4),.w(w10_3),.acc(r10_3),.res(r10_4),.clk(clk),.wout(w10_4));
	PE pe10_5(.x(x5),.w(w10_4),.acc(r10_4),.res(r10_5),.clk(clk),.wout(w10_5));
	PE pe10_6(.x(x6),.w(w10_5),.acc(r10_5),.res(r10_6),.clk(clk),.wout(w10_6));
	PE pe10_7(.x(x7),.w(w10_6),.acc(r10_6),.res(r10_7),.clk(clk),.wout(w10_7));
	PE pe10_8(.x(x8),.w(w10_7),.acc(r10_7),.res(r10_8),.clk(clk),.wout(w10_8));
	PE pe10_9(.x(x9),.w(w10_8),.acc(r10_8),.res(r10_9),.clk(clk),.wout(w10_9));
	PE pe10_10(.x(x10),.w(w10_9),.acc(r10_9),.res(r10_10),.clk(clk),.wout(w10_10));
	PE pe10_11(.x(x11),.w(w10_10),.acc(r10_10),.res(r10_11),.clk(clk),.wout(w10_11));
	PE pe10_12(.x(x12),.w(w10_11),.acc(r10_11),.res(r10_12),.clk(clk),.wout(w10_12));
	PE pe10_13(.x(x13),.w(w10_12),.acc(r10_12),.res(r10_13),.clk(clk),.wout(w10_13));
	PE pe10_14(.x(x14),.w(w10_13),.acc(r10_13),.res(r10_14),.clk(clk),.wout(w10_14));
	PE pe10_15(.x(x15),.w(w10_14),.acc(r10_14),.res(r10_15),.clk(clk),.wout(w10_15));
	PE pe10_16(.x(x16),.w(w10_15),.acc(r10_15),.res(r10_16),.clk(clk),.wout(w10_16));
	PE pe10_17(.x(x17),.w(w10_16),.acc(r10_16),.res(r10_17),.clk(clk),.wout(w10_17));
	PE pe10_18(.x(x18),.w(w10_17),.acc(r10_17),.res(r10_18),.clk(clk),.wout(w10_18));
	PE pe10_19(.x(x19),.w(w10_18),.acc(r10_18),.res(r10_19),.clk(clk),.wout(w10_19));
	PE pe10_20(.x(x20),.w(w10_19),.acc(r10_19),.res(r10_20),.clk(clk),.wout(w10_20));
	PE pe10_21(.x(x21),.w(w10_20),.acc(r10_20),.res(r10_21),.clk(clk),.wout(w10_21));
	PE pe10_22(.x(x22),.w(w10_21),.acc(r10_21),.res(r10_22),.clk(clk),.wout(w10_22));
	PE pe10_23(.x(x23),.w(w10_22),.acc(r10_22),.res(r10_23),.clk(clk),.wout(w10_23));
	PE pe10_24(.x(x24),.w(w10_23),.acc(r10_23),.res(r10_24),.clk(clk),.wout(w10_24));
	PE pe10_25(.x(x25),.w(w10_24),.acc(r10_24),.res(r10_25),.clk(clk),.wout(w10_25));
	PE pe10_26(.x(x26),.w(w10_25),.acc(r10_25),.res(r10_26),.clk(clk),.wout(w10_26));
	PE pe10_27(.x(x27),.w(w10_26),.acc(r10_26),.res(r10_27),.clk(clk),.wout(w10_27));
	PE pe10_28(.x(x28),.w(w10_27),.acc(r10_27),.res(r10_28),.clk(clk),.wout(w10_28));
	PE pe10_29(.x(x29),.w(w10_28),.acc(r10_28),.res(r10_29),.clk(clk),.wout(w10_29));
	PE pe10_30(.x(x30),.w(w10_29),.acc(r10_29),.res(r10_30),.clk(clk),.wout(w10_30));
	PE pe10_31(.x(x31),.w(w10_30),.acc(r10_30),.res(r10_31),.clk(clk),.wout(w10_31));
	PE pe10_32(.x(x32),.w(w10_31),.acc(r10_31),.res(r10_32),.clk(clk),.wout(w10_32));
	PE pe10_33(.x(x33),.w(w10_32),.acc(r10_32),.res(r10_33),.clk(clk),.wout(w10_33));
	PE pe10_34(.x(x34),.w(w10_33),.acc(r10_33),.res(r10_34),.clk(clk),.wout(w10_34));
	PE pe10_35(.x(x35),.w(w10_34),.acc(r10_34),.res(r10_35),.clk(clk),.wout(w10_35));
	PE pe10_36(.x(x36),.w(w10_35),.acc(r10_35),.res(r10_36),.clk(clk),.wout(w10_36));
	PE pe10_37(.x(x37),.w(w10_36),.acc(r10_36),.res(r10_37),.clk(clk),.wout(w10_37));
	PE pe10_38(.x(x38),.w(w10_37),.acc(r10_37),.res(r10_38),.clk(clk),.wout(w10_38));
	PE pe10_39(.x(x39),.w(w10_38),.acc(r10_38),.res(r10_39),.clk(clk),.wout(w10_39));
	PE pe10_40(.x(x40),.w(w10_39),.acc(r10_39),.res(r10_40),.clk(clk),.wout(w10_40));
	PE pe10_41(.x(x41),.w(w10_40),.acc(r10_40),.res(r10_41),.clk(clk),.wout(w10_41));
	PE pe10_42(.x(x42),.w(w10_41),.acc(r10_41),.res(r10_42),.clk(clk),.wout(w10_42));
	PE pe10_43(.x(x43),.w(w10_42),.acc(r10_42),.res(r10_43),.clk(clk),.wout(w10_43));
	PE pe10_44(.x(x44),.w(w10_43),.acc(r10_43),.res(r10_44),.clk(clk),.wout(w10_44));
	PE pe10_45(.x(x45),.w(w10_44),.acc(r10_44),.res(r10_45),.clk(clk),.wout(w10_45));
	PE pe10_46(.x(x46),.w(w10_45),.acc(r10_45),.res(r10_46),.clk(clk),.wout(w10_46));
	PE pe10_47(.x(x47),.w(w10_46),.acc(r10_46),.res(r10_47),.clk(clk),.wout(w10_47));
	PE pe10_48(.x(x48),.w(w10_47),.acc(r10_47),.res(r10_48),.clk(clk),.wout(w10_48));
	PE pe10_49(.x(x49),.w(w10_48),.acc(r10_48),.res(r10_49),.clk(clk),.wout(w10_49));
	PE pe10_50(.x(x50),.w(w10_49),.acc(r10_49),.res(r10_50),.clk(clk),.wout(w10_50));
	PE pe10_51(.x(x51),.w(w10_50),.acc(r10_50),.res(r10_51),.clk(clk),.wout(w10_51));
	PE pe10_52(.x(x52),.w(w10_51),.acc(r10_51),.res(r10_52),.clk(clk),.wout(w10_52));
	PE pe10_53(.x(x53),.w(w10_52),.acc(r10_52),.res(r10_53),.clk(clk),.wout(w10_53));
	PE pe10_54(.x(x54),.w(w10_53),.acc(r10_53),.res(r10_54),.clk(clk),.wout(w10_54));
	PE pe10_55(.x(x55),.w(w10_54),.acc(r10_54),.res(r10_55),.clk(clk),.wout(w10_55));
	PE pe10_56(.x(x56),.w(w10_55),.acc(r10_55),.res(r10_56),.clk(clk),.wout(w10_56));
	PE pe10_57(.x(x57),.w(w10_56),.acc(r10_56),.res(r10_57),.clk(clk),.wout(w10_57));
	PE pe10_58(.x(x58),.w(w10_57),.acc(r10_57),.res(r10_58),.clk(clk),.wout(w10_58));
	PE pe10_59(.x(x59),.w(w10_58),.acc(r10_58),.res(r10_59),.clk(clk),.wout(w10_59));
	PE pe10_60(.x(x60),.w(w10_59),.acc(r10_59),.res(r10_60),.clk(clk),.wout(w10_60));
	PE pe10_61(.x(x61),.w(w10_60),.acc(r10_60),.res(r10_61),.clk(clk),.wout(w10_61));
	PE pe10_62(.x(x62),.w(w10_61),.acc(r10_61),.res(r10_62),.clk(clk),.wout(w10_62));
	PE pe10_63(.x(x63),.w(w10_62),.acc(r10_62),.res(r10_63),.clk(clk),.wout(w10_63));
	PE pe10_64(.x(x64),.w(w10_63),.acc(r10_63),.res(r10_64),.clk(clk),.wout(w10_64));
	PE pe10_65(.x(x65),.w(w10_64),.acc(r10_64),.res(r10_65),.clk(clk),.wout(w10_65));
	PE pe10_66(.x(x66),.w(w10_65),.acc(r10_65),.res(r10_66),.clk(clk),.wout(w10_66));
	PE pe10_67(.x(x67),.w(w10_66),.acc(r10_66),.res(r10_67),.clk(clk),.wout(w10_67));
	PE pe10_68(.x(x68),.w(w10_67),.acc(r10_67),.res(r10_68),.clk(clk),.wout(w10_68));
	PE pe10_69(.x(x69),.w(w10_68),.acc(r10_68),.res(r10_69),.clk(clk),.wout(w10_69));
	PE pe10_70(.x(x70),.w(w10_69),.acc(r10_69),.res(r10_70),.clk(clk),.wout(w10_70));
	PE pe10_71(.x(x71),.w(w10_70),.acc(r10_70),.res(r10_71),.clk(clk),.wout(w10_71));
	PE pe10_72(.x(x72),.w(w10_71),.acc(r10_71),.res(r10_72),.clk(clk),.wout(w10_72));
	PE pe10_73(.x(x73),.w(w10_72),.acc(r10_72),.res(r10_73),.clk(clk),.wout(w10_73));
	PE pe10_74(.x(x74),.w(w10_73),.acc(r10_73),.res(r10_74),.clk(clk),.wout(w10_74));
	PE pe10_75(.x(x75),.w(w10_74),.acc(r10_74),.res(r10_75),.clk(clk),.wout(w10_75));
	PE pe10_76(.x(x76),.w(w10_75),.acc(r10_75),.res(r10_76),.clk(clk),.wout(w10_76));
	PE pe10_77(.x(x77),.w(w10_76),.acc(r10_76),.res(r10_77),.clk(clk),.wout(w10_77));
	PE pe10_78(.x(x78),.w(w10_77),.acc(r10_77),.res(r10_78),.clk(clk),.wout(w10_78));
	PE pe10_79(.x(x79),.w(w10_78),.acc(r10_78),.res(r10_79),.clk(clk),.wout(w10_79));
	PE pe10_80(.x(x80),.w(w10_79),.acc(r10_79),.res(r10_80),.clk(clk),.wout(w10_80));
	PE pe10_81(.x(x81),.w(w10_80),.acc(r10_80),.res(r10_81),.clk(clk),.wout(w10_81));
	PE pe10_82(.x(x82),.w(w10_81),.acc(r10_81),.res(r10_82),.clk(clk),.wout(w10_82));
	PE pe10_83(.x(x83),.w(w10_82),.acc(r10_82),.res(r10_83),.clk(clk),.wout(w10_83));
	PE pe10_84(.x(x84),.w(w10_83),.acc(r10_83),.res(r10_84),.clk(clk),.wout(w10_84));
	PE pe10_85(.x(x85),.w(w10_84),.acc(r10_84),.res(r10_85),.clk(clk),.wout(w10_85));
	PE pe10_86(.x(x86),.w(w10_85),.acc(r10_85),.res(r10_86),.clk(clk),.wout(w10_86));
	PE pe10_87(.x(x87),.w(w10_86),.acc(r10_86),.res(r10_87),.clk(clk),.wout(w10_87));
	PE pe10_88(.x(x88),.w(w10_87),.acc(r10_87),.res(r10_88),.clk(clk),.wout(w10_88));
	PE pe10_89(.x(x89),.w(w10_88),.acc(r10_88),.res(r10_89),.clk(clk),.wout(w10_89));
	PE pe10_90(.x(x90),.w(w10_89),.acc(r10_89),.res(r10_90),.clk(clk),.wout(w10_90));
	PE pe10_91(.x(x91),.w(w10_90),.acc(r10_90),.res(r10_91),.clk(clk),.wout(w10_91));
	PE pe10_92(.x(x92),.w(w10_91),.acc(r10_91),.res(r10_92),.clk(clk),.wout(w10_92));
	PE pe10_93(.x(x93),.w(w10_92),.acc(r10_92),.res(r10_93),.clk(clk),.wout(w10_93));
	PE pe10_94(.x(x94),.w(w10_93),.acc(r10_93),.res(r10_94),.clk(clk),.wout(w10_94));
	PE pe10_95(.x(x95),.w(w10_94),.acc(r10_94),.res(r10_95),.clk(clk),.wout(w10_95));
	PE pe10_96(.x(x96),.w(w10_95),.acc(r10_95),.res(r10_96),.clk(clk),.wout(w10_96));
	PE pe10_97(.x(x97),.w(w10_96),.acc(r10_96),.res(r10_97),.clk(clk),.wout(w10_97));
	PE pe10_98(.x(x98),.w(w10_97),.acc(r10_97),.res(r10_98),.clk(clk),.wout(w10_98));
	PE pe10_99(.x(x99),.w(w10_98),.acc(r10_98),.res(r10_99),.clk(clk),.wout(w10_99));
	PE pe10_100(.x(x100),.w(w10_99),.acc(r10_99),.res(r10_100),.clk(clk),.wout(w10_100));
	PE pe10_101(.x(x101),.w(w10_100),.acc(r10_100),.res(r10_101),.clk(clk),.wout(w10_101));
	PE pe10_102(.x(x102),.w(w10_101),.acc(r10_101),.res(r10_102),.clk(clk),.wout(w10_102));
	PE pe10_103(.x(x103),.w(w10_102),.acc(r10_102),.res(r10_103),.clk(clk),.wout(w10_103));
	PE pe10_104(.x(x104),.w(w10_103),.acc(r10_103),.res(r10_104),.clk(clk),.wout(w10_104));
	PE pe10_105(.x(x105),.w(w10_104),.acc(r10_104),.res(r10_105),.clk(clk),.wout(w10_105));
	PE pe10_106(.x(x106),.w(w10_105),.acc(r10_105),.res(r10_106),.clk(clk),.wout(w10_106));
	PE pe10_107(.x(x107),.w(w10_106),.acc(r10_106),.res(r10_107),.clk(clk),.wout(w10_107));
	PE pe10_108(.x(x108),.w(w10_107),.acc(r10_107),.res(r10_108),.clk(clk),.wout(w10_108));
	PE pe10_109(.x(x109),.w(w10_108),.acc(r10_108),.res(r10_109),.clk(clk),.wout(w10_109));
	PE pe10_110(.x(x110),.w(w10_109),.acc(r10_109),.res(r10_110),.clk(clk),.wout(w10_110));
	PE pe10_111(.x(x111),.w(w10_110),.acc(r10_110),.res(r10_111),.clk(clk),.wout(w10_111));
	PE pe10_112(.x(x112),.w(w10_111),.acc(r10_111),.res(r10_112),.clk(clk),.wout(w10_112));
	PE pe10_113(.x(x113),.w(w10_112),.acc(r10_112),.res(r10_113),.clk(clk),.wout(w10_113));
	PE pe10_114(.x(x114),.w(w10_113),.acc(r10_113),.res(r10_114),.clk(clk),.wout(w10_114));
	PE pe10_115(.x(x115),.w(w10_114),.acc(r10_114),.res(r10_115),.clk(clk),.wout(w10_115));
	PE pe10_116(.x(x116),.w(w10_115),.acc(r10_115),.res(r10_116),.clk(clk),.wout(w10_116));
	PE pe10_117(.x(x117),.w(w10_116),.acc(r10_116),.res(r10_117),.clk(clk),.wout(w10_117));
	PE pe10_118(.x(x118),.w(w10_117),.acc(r10_117),.res(r10_118),.clk(clk),.wout(w10_118));
	PE pe10_119(.x(x119),.w(w10_118),.acc(r10_118),.res(r10_119),.clk(clk),.wout(w10_119));
	PE pe10_120(.x(x120),.w(w10_119),.acc(r10_119),.res(r10_120),.clk(clk),.wout(w10_120));
	PE pe10_121(.x(x121),.w(w10_120),.acc(r10_120),.res(r10_121),.clk(clk),.wout(w10_121));
	PE pe10_122(.x(x122),.w(w10_121),.acc(r10_121),.res(r10_122),.clk(clk),.wout(w10_122));
	PE pe10_123(.x(x123),.w(w10_122),.acc(r10_122),.res(r10_123),.clk(clk),.wout(w10_123));
	PE pe10_124(.x(x124),.w(w10_123),.acc(r10_123),.res(r10_124),.clk(clk),.wout(w10_124));
	PE pe10_125(.x(x125),.w(w10_124),.acc(r10_124),.res(r10_125),.clk(clk),.wout(w10_125));
	PE pe10_126(.x(x126),.w(w10_125),.acc(r10_125),.res(r10_126),.clk(clk),.wout(w10_126));
	PE pe10_127(.x(x127),.w(w10_126),.acc(r10_126),.res(result10),.clk(clk),.wout(weight10));

	PE pe11_0(.x(x0),.w(w11),.acc(32'h0),.res(r11_0),.clk(clk),.wout(w11_0));
	PE pe11_1(.x(x1),.w(w11_0),.acc(r11_0),.res(r11_1),.clk(clk),.wout(w11_1));
	PE pe11_2(.x(x2),.w(w11_1),.acc(r11_1),.res(r11_2),.clk(clk),.wout(w11_2));
	PE pe11_3(.x(x3),.w(w11_2),.acc(r11_2),.res(r11_3),.clk(clk),.wout(w11_3));
	PE pe11_4(.x(x4),.w(w11_3),.acc(r11_3),.res(r11_4),.clk(clk),.wout(w11_4));
	PE pe11_5(.x(x5),.w(w11_4),.acc(r11_4),.res(r11_5),.clk(clk),.wout(w11_5));
	PE pe11_6(.x(x6),.w(w11_5),.acc(r11_5),.res(r11_6),.clk(clk),.wout(w11_6));
	PE pe11_7(.x(x7),.w(w11_6),.acc(r11_6),.res(r11_7),.clk(clk),.wout(w11_7));
	PE pe11_8(.x(x8),.w(w11_7),.acc(r11_7),.res(r11_8),.clk(clk),.wout(w11_8));
	PE pe11_9(.x(x9),.w(w11_8),.acc(r11_8),.res(r11_9),.clk(clk),.wout(w11_9));
	PE pe11_10(.x(x10),.w(w11_9),.acc(r11_9),.res(r11_10),.clk(clk),.wout(w11_10));
	PE pe11_11(.x(x11),.w(w11_10),.acc(r11_10),.res(r11_11),.clk(clk),.wout(w11_11));
	PE pe11_12(.x(x12),.w(w11_11),.acc(r11_11),.res(r11_12),.clk(clk),.wout(w11_12));
	PE pe11_13(.x(x13),.w(w11_12),.acc(r11_12),.res(r11_13),.clk(clk),.wout(w11_13));
	PE pe11_14(.x(x14),.w(w11_13),.acc(r11_13),.res(r11_14),.clk(clk),.wout(w11_14));
	PE pe11_15(.x(x15),.w(w11_14),.acc(r11_14),.res(r11_15),.clk(clk),.wout(w11_15));
	PE pe11_16(.x(x16),.w(w11_15),.acc(r11_15),.res(r11_16),.clk(clk),.wout(w11_16));
	PE pe11_17(.x(x17),.w(w11_16),.acc(r11_16),.res(r11_17),.clk(clk),.wout(w11_17));
	PE pe11_18(.x(x18),.w(w11_17),.acc(r11_17),.res(r11_18),.clk(clk),.wout(w11_18));
	PE pe11_19(.x(x19),.w(w11_18),.acc(r11_18),.res(r11_19),.clk(clk),.wout(w11_19));
	PE pe11_20(.x(x20),.w(w11_19),.acc(r11_19),.res(r11_20),.clk(clk),.wout(w11_20));
	PE pe11_21(.x(x21),.w(w11_20),.acc(r11_20),.res(r11_21),.clk(clk),.wout(w11_21));
	PE pe11_22(.x(x22),.w(w11_21),.acc(r11_21),.res(r11_22),.clk(clk),.wout(w11_22));
	PE pe11_23(.x(x23),.w(w11_22),.acc(r11_22),.res(r11_23),.clk(clk),.wout(w11_23));
	PE pe11_24(.x(x24),.w(w11_23),.acc(r11_23),.res(r11_24),.clk(clk),.wout(w11_24));
	PE pe11_25(.x(x25),.w(w11_24),.acc(r11_24),.res(r11_25),.clk(clk),.wout(w11_25));
	PE pe11_26(.x(x26),.w(w11_25),.acc(r11_25),.res(r11_26),.clk(clk),.wout(w11_26));
	PE pe11_27(.x(x27),.w(w11_26),.acc(r11_26),.res(r11_27),.clk(clk),.wout(w11_27));
	PE pe11_28(.x(x28),.w(w11_27),.acc(r11_27),.res(r11_28),.clk(clk),.wout(w11_28));
	PE pe11_29(.x(x29),.w(w11_28),.acc(r11_28),.res(r11_29),.clk(clk),.wout(w11_29));
	PE pe11_30(.x(x30),.w(w11_29),.acc(r11_29),.res(r11_30),.clk(clk),.wout(w11_30));
	PE pe11_31(.x(x31),.w(w11_30),.acc(r11_30),.res(r11_31),.clk(clk),.wout(w11_31));
	PE pe11_32(.x(x32),.w(w11_31),.acc(r11_31),.res(r11_32),.clk(clk),.wout(w11_32));
	PE pe11_33(.x(x33),.w(w11_32),.acc(r11_32),.res(r11_33),.clk(clk),.wout(w11_33));
	PE pe11_34(.x(x34),.w(w11_33),.acc(r11_33),.res(r11_34),.clk(clk),.wout(w11_34));
	PE pe11_35(.x(x35),.w(w11_34),.acc(r11_34),.res(r11_35),.clk(clk),.wout(w11_35));
	PE pe11_36(.x(x36),.w(w11_35),.acc(r11_35),.res(r11_36),.clk(clk),.wout(w11_36));
	PE pe11_37(.x(x37),.w(w11_36),.acc(r11_36),.res(r11_37),.clk(clk),.wout(w11_37));
	PE pe11_38(.x(x38),.w(w11_37),.acc(r11_37),.res(r11_38),.clk(clk),.wout(w11_38));
	PE pe11_39(.x(x39),.w(w11_38),.acc(r11_38),.res(r11_39),.clk(clk),.wout(w11_39));
	PE pe11_40(.x(x40),.w(w11_39),.acc(r11_39),.res(r11_40),.clk(clk),.wout(w11_40));
	PE pe11_41(.x(x41),.w(w11_40),.acc(r11_40),.res(r11_41),.clk(clk),.wout(w11_41));
	PE pe11_42(.x(x42),.w(w11_41),.acc(r11_41),.res(r11_42),.clk(clk),.wout(w11_42));
	PE pe11_43(.x(x43),.w(w11_42),.acc(r11_42),.res(r11_43),.clk(clk),.wout(w11_43));
	PE pe11_44(.x(x44),.w(w11_43),.acc(r11_43),.res(r11_44),.clk(clk),.wout(w11_44));
	PE pe11_45(.x(x45),.w(w11_44),.acc(r11_44),.res(r11_45),.clk(clk),.wout(w11_45));
	PE pe11_46(.x(x46),.w(w11_45),.acc(r11_45),.res(r11_46),.clk(clk),.wout(w11_46));
	PE pe11_47(.x(x47),.w(w11_46),.acc(r11_46),.res(r11_47),.clk(clk),.wout(w11_47));
	PE pe11_48(.x(x48),.w(w11_47),.acc(r11_47),.res(r11_48),.clk(clk),.wout(w11_48));
	PE pe11_49(.x(x49),.w(w11_48),.acc(r11_48),.res(r11_49),.clk(clk),.wout(w11_49));
	PE pe11_50(.x(x50),.w(w11_49),.acc(r11_49),.res(r11_50),.clk(clk),.wout(w11_50));
	PE pe11_51(.x(x51),.w(w11_50),.acc(r11_50),.res(r11_51),.clk(clk),.wout(w11_51));
	PE pe11_52(.x(x52),.w(w11_51),.acc(r11_51),.res(r11_52),.clk(clk),.wout(w11_52));
	PE pe11_53(.x(x53),.w(w11_52),.acc(r11_52),.res(r11_53),.clk(clk),.wout(w11_53));
	PE pe11_54(.x(x54),.w(w11_53),.acc(r11_53),.res(r11_54),.clk(clk),.wout(w11_54));
	PE pe11_55(.x(x55),.w(w11_54),.acc(r11_54),.res(r11_55),.clk(clk),.wout(w11_55));
	PE pe11_56(.x(x56),.w(w11_55),.acc(r11_55),.res(r11_56),.clk(clk),.wout(w11_56));
	PE pe11_57(.x(x57),.w(w11_56),.acc(r11_56),.res(r11_57),.clk(clk),.wout(w11_57));
	PE pe11_58(.x(x58),.w(w11_57),.acc(r11_57),.res(r11_58),.clk(clk),.wout(w11_58));
	PE pe11_59(.x(x59),.w(w11_58),.acc(r11_58),.res(r11_59),.clk(clk),.wout(w11_59));
	PE pe11_60(.x(x60),.w(w11_59),.acc(r11_59),.res(r11_60),.clk(clk),.wout(w11_60));
	PE pe11_61(.x(x61),.w(w11_60),.acc(r11_60),.res(r11_61),.clk(clk),.wout(w11_61));
	PE pe11_62(.x(x62),.w(w11_61),.acc(r11_61),.res(r11_62),.clk(clk),.wout(w11_62));
	PE pe11_63(.x(x63),.w(w11_62),.acc(r11_62),.res(r11_63),.clk(clk),.wout(w11_63));
	PE pe11_64(.x(x64),.w(w11_63),.acc(r11_63),.res(r11_64),.clk(clk),.wout(w11_64));
	PE pe11_65(.x(x65),.w(w11_64),.acc(r11_64),.res(r11_65),.clk(clk),.wout(w11_65));
	PE pe11_66(.x(x66),.w(w11_65),.acc(r11_65),.res(r11_66),.clk(clk),.wout(w11_66));
	PE pe11_67(.x(x67),.w(w11_66),.acc(r11_66),.res(r11_67),.clk(clk),.wout(w11_67));
	PE pe11_68(.x(x68),.w(w11_67),.acc(r11_67),.res(r11_68),.clk(clk),.wout(w11_68));
	PE pe11_69(.x(x69),.w(w11_68),.acc(r11_68),.res(r11_69),.clk(clk),.wout(w11_69));
	PE pe11_70(.x(x70),.w(w11_69),.acc(r11_69),.res(r11_70),.clk(clk),.wout(w11_70));
	PE pe11_71(.x(x71),.w(w11_70),.acc(r11_70),.res(r11_71),.clk(clk),.wout(w11_71));
	PE pe11_72(.x(x72),.w(w11_71),.acc(r11_71),.res(r11_72),.clk(clk),.wout(w11_72));
	PE pe11_73(.x(x73),.w(w11_72),.acc(r11_72),.res(r11_73),.clk(clk),.wout(w11_73));
	PE pe11_74(.x(x74),.w(w11_73),.acc(r11_73),.res(r11_74),.clk(clk),.wout(w11_74));
	PE pe11_75(.x(x75),.w(w11_74),.acc(r11_74),.res(r11_75),.clk(clk),.wout(w11_75));
	PE pe11_76(.x(x76),.w(w11_75),.acc(r11_75),.res(r11_76),.clk(clk),.wout(w11_76));
	PE pe11_77(.x(x77),.w(w11_76),.acc(r11_76),.res(r11_77),.clk(clk),.wout(w11_77));
	PE pe11_78(.x(x78),.w(w11_77),.acc(r11_77),.res(r11_78),.clk(clk),.wout(w11_78));
	PE pe11_79(.x(x79),.w(w11_78),.acc(r11_78),.res(r11_79),.clk(clk),.wout(w11_79));
	PE pe11_80(.x(x80),.w(w11_79),.acc(r11_79),.res(r11_80),.clk(clk),.wout(w11_80));
	PE pe11_81(.x(x81),.w(w11_80),.acc(r11_80),.res(r11_81),.clk(clk),.wout(w11_81));
	PE pe11_82(.x(x82),.w(w11_81),.acc(r11_81),.res(r11_82),.clk(clk),.wout(w11_82));
	PE pe11_83(.x(x83),.w(w11_82),.acc(r11_82),.res(r11_83),.clk(clk),.wout(w11_83));
	PE pe11_84(.x(x84),.w(w11_83),.acc(r11_83),.res(r11_84),.clk(clk),.wout(w11_84));
	PE pe11_85(.x(x85),.w(w11_84),.acc(r11_84),.res(r11_85),.clk(clk),.wout(w11_85));
	PE pe11_86(.x(x86),.w(w11_85),.acc(r11_85),.res(r11_86),.clk(clk),.wout(w11_86));
	PE pe11_87(.x(x87),.w(w11_86),.acc(r11_86),.res(r11_87),.clk(clk),.wout(w11_87));
	PE pe11_88(.x(x88),.w(w11_87),.acc(r11_87),.res(r11_88),.clk(clk),.wout(w11_88));
	PE pe11_89(.x(x89),.w(w11_88),.acc(r11_88),.res(r11_89),.clk(clk),.wout(w11_89));
	PE pe11_90(.x(x90),.w(w11_89),.acc(r11_89),.res(r11_90),.clk(clk),.wout(w11_90));
	PE pe11_91(.x(x91),.w(w11_90),.acc(r11_90),.res(r11_91),.clk(clk),.wout(w11_91));
	PE pe11_92(.x(x92),.w(w11_91),.acc(r11_91),.res(r11_92),.clk(clk),.wout(w11_92));
	PE pe11_93(.x(x93),.w(w11_92),.acc(r11_92),.res(r11_93),.clk(clk),.wout(w11_93));
	PE pe11_94(.x(x94),.w(w11_93),.acc(r11_93),.res(r11_94),.clk(clk),.wout(w11_94));
	PE pe11_95(.x(x95),.w(w11_94),.acc(r11_94),.res(r11_95),.clk(clk),.wout(w11_95));
	PE pe11_96(.x(x96),.w(w11_95),.acc(r11_95),.res(r11_96),.clk(clk),.wout(w11_96));
	PE pe11_97(.x(x97),.w(w11_96),.acc(r11_96),.res(r11_97),.clk(clk),.wout(w11_97));
	PE pe11_98(.x(x98),.w(w11_97),.acc(r11_97),.res(r11_98),.clk(clk),.wout(w11_98));
	PE pe11_99(.x(x99),.w(w11_98),.acc(r11_98),.res(r11_99),.clk(clk),.wout(w11_99));
	PE pe11_100(.x(x100),.w(w11_99),.acc(r11_99),.res(r11_100),.clk(clk),.wout(w11_100));
	PE pe11_101(.x(x101),.w(w11_100),.acc(r11_100),.res(r11_101),.clk(clk),.wout(w11_101));
	PE pe11_102(.x(x102),.w(w11_101),.acc(r11_101),.res(r11_102),.clk(clk),.wout(w11_102));
	PE pe11_103(.x(x103),.w(w11_102),.acc(r11_102),.res(r11_103),.clk(clk),.wout(w11_103));
	PE pe11_104(.x(x104),.w(w11_103),.acc(r11_103),.res(r11_104),.clk(clk),.wout(w11_104));
	PE pe11_105(.x(x105),.w(w11_104),.acc(r11_104),.res(r11_105),.clk(clk),.wout(w11_105));
	PE pe11_106(.x(x106),.w(w11_105),.acc(r11_105),.res(r11_106),.clk(clk),.wout(w11_106));
	PE pe11_107(.x(x107),.w(w11_106),.acc(r11_106),.res(r11_107),.clk(clk),.wout(w11_107));
	PE pe11_108(.x(x108),.w(w11_107),.acc(r11_107),.res(r11_108),.clk(clk),.wout(w11_108));
	PE pe11_109(.x(x109),.w(w11_108),.acc(r11_108),.res(r11_109),.clk(clk),.wout(w11_109));
	PE pe11_110(.x(x110),.w(w11_109),.acc(r11_109),.res(r11_110),.clk(clk),.wout(w11_110));
	PE pe11_111(.x(x111),.w(w11_110),.acc(r11_110),.res(r11_111),.clk(clk),.wout(w11_111));
	PE pe11_112(.x(x112),.w(w11_111),.acc(r11_111),.res(r11_112),.clk(clk),.wout(w11_112));
	PE pe11_113(.x(x113),.w(w11_112),.acc(r11_112),.res(r11_113),.clk(clk),.wout(w11_113));
	PE pe11_114(.x(x114),.w(w11_113),.acc(r11_113),.res(r11_114),.clk(clk),.wout(w11_114));
	PE pe11_115(.x(x115),.w(w11_114),.acc(r11_114),.res(r11_115),.clk(clk),.wout(w11_115));
	PE pe11_116(.x(x116),.w(w11_115),.acc(r11_115),.res(r11_116),.clk(clk),.wout(w11_116));
	PE pe11_117(.x(x117),.w(w11_116),.acc(r11_116),.res(r11_117),.clk(clk),.wout(w11_117));
	PE pe11_118(.x(x118),.w(w11_117),.acc(r11_117),.res(r11_118),.clk(clk),.wout(w11_118));
	PE pe11_119(.x(x119),.w(w11_118),.acc(r11_118),.res(r11_119),.clk(clk),.wout(w11_119));
	PE pe11_120(.x(x120),.w(w11_119),.acc(r11_119),.res(r11_120),.clk(clk),.wout(w11_120));
	PE pe11_121(.x(x121),.w(w11_120),.acc(r11_120),.res(r11_121),.clk(clk),.wout(w11_121));
	PE pe11_122(.x(x122),.w(w11_121),.acc(r11_121),.res(r11_122),.clk(clk),.wout(w11_122));
	PE pe11_123(.x(x123),.w(w11_122),.acc(r11_122),.res(r11_123),.clk(clk),.wout(w11_123));
	PE pe11_124(.x(x124),.w(w11_123),.acc(r11_123),.res(r11_124),.clk(clk),.wout(w11_124));
	PE pe11_125(.x(x125),.w(w11_124),.acc(r11_124),.res(r11_125),.clk(clk),.wout(w11_125));
	PE pe11_126(.x(x126),.w(w11_125),.acc(r11_125),.res(r11_126),.clk(clk),.wout(w11_126));
	PE pe11_127(.x(x127),.w(w11_126),.acc(r11_126),.res(result11),.clk(clk),.wout(weight11));

	PE pe12_0(.x(x0),.w(w12),.acc(32'h0),.res(r12_0),.clk(clk),.wout(w12_0));
	PE pe12_1(.x(x1),.w(w12_0),.acc(r12_0),.res(r12_1),.clk(clk),.wout(w12_1));
	PE pe12_2(.x(x2),.w(w12_1),.acc(r12_1),.res(r12_2),.clk(clk),.wout(w12_2));
	PE pe12_3(.x(x3),.w(w12_2),.acc(r12_2),.res(r12_3),.clk(clk),.wout(w12_3));
	PE pe12_4(.x(x4),.w(w12_3),.acc(r12_3),.res(r12_4),.clk(clk),.wout(w12_4));
	PE pe12_5(.x(x5),.w(w12_4),.acc(r12_4),.res(r12_5),.clk(clk),.wout(w12_5));
	PE pe12_6(.x(x6),.w(w12_5),.acc(r12_5),.res(r12_6),.clk(clk),.wout(w12_6));
	PE pe12_7(.x(x7),.w(w12_6),.acc(r12_6),.res(r12_7),.clk(clk),.wout(w12_7));
	PE pe12_8(.x(x8),.w(w12_7),.acc(r12_7),.res(r12_8),.clk(clk),.wout(w12_8));
	PE pe12_9(.x(x9),.w(w12_8),.acc(r12_8),.res(r12_9),.clk(clk),.wout(w12_9));
	PE pe12_10(.x(x10),.w(w12_9),.acc(r12_9),.res(r12_10),.clk(clk),.wout(w12_10));
	PE pe12_11(.x(x11),.w(w12_10),.acc(r12_10),.res(r12_11),.clk(clk),.wout(w12_11));
	PE pe12_12(.x(x12),.w(w12_11),.acc(r12_11),.res(r12_12),.clk(clk),.wout(w12_12));
	PE pe12_13(.x(x13),.w(w12_12),.acc(r12_12),.res(r12_13),.clk(clk),.wout(w12_13));
	PE pe12_14(.x(x14),.w(w12_13),.acc(r12_13),.res(r12_14),.clk(clk),.wout(w12_14));
	PE pe12_15(.x(x15),.w(w12_14),.acc(r12_14),.res(r12_15),.clk(clk),.wout(w12_15));
	PE pe12_16(.x(x16),.w(w12_15),.acc(r12_15),.res(r12_16),.clk(clk),.wout(w12_16));
	PE pe12_17(.x(x17),.w(w12_16),.acc(r12_16),.res(r12_17),.clk(clk),.wout(w12_17));
	PE pe12_18(.x(x18),.w(w12_17),.acc(r12_17),.res(r12_18),.clk(clk),.wout(w12_18));
	PE pe12_19(.x(x19),.w(w12_18),.acc(r12_18),.res(r12_19),.clk(clk),.wout(w12_19));
	PE pe12_20(.x(x20),.w(w12_19),.acc(r12_19),.res(r12_20),.clk(clk),.wout(w12_20));
	PE pe12_21(.x(x21),.w(w12_20),.acc(r12_20),.res(r12_21),.clk(clk),.wout(w12_21));
	PE pe12_22(.x(x22),.w(w12_21),.acc(r12_21),.res(r12_22),.clk(clk),.wout(w12_22));
	PE pe12_23(.x(x23),.w(w12_22),.acc(r12_22),.res(r12_23),.clk(clk),.wout(w12_23));
	PE pe12_24(.x(x24),.w(w12_23),.acc(r12_23),.res(r12_24),.clk(clk),.wout(w12_24));
	PE pe12_25(.x(x25),.w(w12_24),.acc(r12_24),.res(r12_25),.clk(clk),.wout(w12_25));
	PE pe12_26(.x(x26),.w(w12_25),.acc(r12_25),.res(r12_26),.clk(clk),.wout(w12_26));
	PE pe12_27(.x(x27),.w(w12_26),.acc(r12_26),.res(r12_27),.clk(clk),.wout(w12_27));
	PE pe12_28(.x(x28),.w(w12_27),.acc(r12_27),.res(r12_28),.clk(clk),.wout(w12_28));
	PE pe12_29(.x(x29),.w(w12_28),.acc(r12_28),.res(r12_29),.clk(clk),.wout(w12_29));
	PE pe12_30(.x(x30),.w(w12_29),.acc(r12_29),.res(r12_30),.clk(clk),.wout(w12_30));
	PE pe12_31(.x(x31),.w(w12_30),.acc(r12_30),.res(r12_31),.clk(clk),.wout(w12_31));
	PE pe12_32(.x(x32),.w(w12_31),.acc(r12_31),.res(r12_32),.clk(clk),.wout(w12_32));
	PE pe12_33(.x(x33),.w(w12_32),.acc(r12_32),.res(r12_33),.clk(clk),.wout(w12_33));
	PE pe12_34(.x(x34),.w(w12_33),.acc(r12_33),.res(r12_34),.clk(clk),.wout(w12_34));
	PE pe12_35(.x(x35),.w(w12_34),.acc(r12_34),.res(r12_35),.clk(clk),.wout(w12_35));
	PE pe12_36(.x(x36),.w(w12_35),.acc(r12_35),.res(r12_36),.clk(clk),.wout(w12_36));
	PE pe12_37(.x(x37),.w(w12_36),.acc(r12_36),.res(r12_37),.clk(clk),.wout(w12_37));
	PE pe12_38(.x(x38),.w(w12_37),.acc(r12_37),.res(r12_38),.clk(clk),.wout(w12_38));
	PE pe12_39(.x(x39),.w(w12_38),.acc(r12_38),.res(r12_39),.clk(clk),.wout(w12_39));
	PE pe12_40(.x(x40),.w(w12_39),.acc(r12_39),.res(r12_40),.clk(clk),.wout(w12_40));
	PE pe12_41(.x(x41),.w(w12_40),.acc(r12_40),.res(r12_41),.clk(clk),.wout(w12_41));
	PE pe12_42(.x(x42),.w(w12_41),.acc(r12_41),.res(r12_42),.clk(clk),.wout(w12_42));
	PE pe12_43(.x(x43),.w(w12_42),.acc(r12_42),.res(r12_43),.clk(clk),.wout(w12_43));
	PE pe12_44(.x(x44),.w(w12_43),.acc(r12_43),.res(r12_44),.clk(clk),.wout(w12_44));
	PE pe12_45(.x(x45),.w(w12_44),.acc(r12_44),.res(r12_45),.clk(clk),.wout(w12_45));
	PE pe12_46(.x(x46),.w(w12_45),.acc(r12_45),.res(r12_46),.clk(clk),.wout(w12_46));
	PE pe12_47(.x(x47),.w(w12_46),.acc(r12_46),.res(r12_47),.clk(clk),.wout(w12_47));
	PE pe12_48(.x(x48),.w(w12_47),.acc(r12_47),.res(r12_48),.clk(clk),.wout(w12_48));
	PE pe12_49(.x(x49),.w(w12_48),.acc(r12_48),.res(r12_49),.clk(clk),.wout(w12_49));
	PE pe12_50(.x(x50),.w(w12_49),.acc(r12_49),.res(r12_50),.clk(clk),.wout(w12_50));
	PE pe12_51(.x(x51),.w(w12_50),.acc(r12_50),.res(r12_51),.clk(clk),.wout(w12_51));
	PE pe12_52(.x(x52),.w(w12_51),.acc(r12_51),.res(r12_52),.clk(clk),.wout(w12_52));
	PE pe12_53(.x(x53),.w(w12_52),.acc(r12_52),.res(r12_53),.clk(clk),.wout(w12_53));
	PE pe12_54(.x(x54),.w(w12_53),.acc(r12_53),.res(r12_54),.clk(clk),.wout(w12_54));
	PE pe12_55(.x(x55),.w(w12_54),.acc(r12_54),.res(r12_55),.clk(clk),.wout(w12_55));
	PE pe12_56(.x(x56),.w(w12_55),.acc(r12_55),.res(r12_56),.clk(clk),.wout(w12_56));
	PE pe12_57(.x(x57),.w(w12_56),.acc(r12_56),.res(r12_57),.clk(clk),.wout(w12_57));
	PE pe12_58(.x(x58),.w(w12_57),.acc(r12_57),.res(r12_58),.clk(clk),.wout(w12_58));
	PE pe12_59(.x(x59),.w(w12_58),.acc(r12_58),.res(r12_59),.clk(clk),.wout(w12_59));
	PE pe12_60(.x(x60),.w(w12_59),.acc(r12_59),.res(r12_60),.clk(clk),.wout(w12_60));
	PE pe12_61(.x(x61),.w(w12_60),.acc(r12_60),.res(r12_61),.clk(clk),.wout(w12_61));
	PE pe12_62(.x(x62),.w(w12_61),.acc(r12_61),.res(r12_62),.clk(clk),.wout(w12_62));
	PE pe12_63(.x(x63),.w(w12_62),.acc(r12_62),.res(r12_63),.clk(clk),.wout(w12_63));
	PE pe12_64(.x(x64),.w(w12_63),.acc(r12_63),.res(r12_64),.clk(clk),.wout(w12_64));
	PE pe12_65(.x(x65),.w(w12_64),.acc(r12_64),.res(r12_65),.clk(clk),.wout(w12_65));
	PE pe12_66(.x(x66),.w(w12_65),.acc(r12_65),.res(r12_66),.clk(clk),.wout(w12_66));
	PE pe12_67(.x(x67),.w(w12_66),.acc(r12_66),.res(r12_67),.clk(clk),.wout(w12_67));
	PE pe12_68(.x(x68),.w(w12_67),.acc(r12_67),.res(r12_68),.clk(clk),.wout(w12_68));
	PE pe12_69(.x(x69),.w(w12_68),.acc(r12_68),.res(r12_69),.clk(clk),.wout(w12_69));
	PE pe12_70(.x(x70),.w(w12_69),.acc(r12_69),.res(r12_70),.clk(clk),.wout(w12_70));
	PE pe12_71(.x(x71),.w(w12_70),.acc(r12_70),.res(r12_71),.clk(clk),.wout(w12_71));
	PE pe12_72(.x(x72),.w(w12_71),.acc(r12_71),.res(r12_72),.clk(clk),.wout(w12_72));
	PE pe12_73(.x(x73),.w(w12_72),.acc(r12_72),.res(r12_73),.clk(clk),.wout(w12_73));
	PE pe12_74(.x(x74),.w(w12_73),.acc(r12_73),.res(r12_74),.clk(clk),.wout(w12_74));
	PE pe12_75(.x(x75),.w(w12_74),.acc(r12_74),.res(r12_75),.clk(clk),.wout(w12_75));
	PE pe12_76(.x(x76),.w(w12_75),.acc(r12_75),.res(r12_76),.clk(clk),.wout(w12_76));
	PE pe12_77(.x(x77),.w(w12_76),.acc(r12_76),.res(r12_77),.clk(clk),.wout(w12_77));
	PE pe12_78(.x(x78),.w(w12_77),.acc(r12_77),.res(r12_78),.clk(clk),.wout(w12_78));
	PE pe12_79(.x(x79),.w(w12_78),.acc(r12_78),.res(r12_79),.clk(clk),.wout(w12_79));
	PE pe12_80(.x(x80),.w(w12_79),.acc(r12_79),.res(r12_80),.clk(clk),.wout(w12_80));
	PE pe12_81(.x(x81),.w(w12_80),.acc(r12_80),.res(r12_81),.clk(clk),.wout(w12_81));
	PE pe12_82(.x(x82),.w(w12_81),.acc(r12_81),.res(r12_82),.clk(clk),.wout(w12_82));
	PE pe12_83(.x(x83),.w(w12_82),.acc(r12_82),.res(r12_83),.clk(clk),.wout(w12_83));
	PE pe12_84(.x(x84),.w(w12_83),.acc(r12_83),.res(r12_84),.clk(clk),.wout(w12_84));
	PE pe12_85(.x(x85),.w(w12_84),.acc(r12_84),.res(r12_85),.clk(clk),.wout(w12_85));
	PE pe12_86(.x(x86),.w(w12_85),.acc(r12_85),.res(r12_86),.clk(clk),.wout(w12_86));
	PE pe12_87(.x(x87),.w(w12_86),.acc(r12_86),.res(r12_87),.clk(clk),.wout(w12_87));
	PE pe12_88(.x(x88),.w(w12_87),.acc(r12_87),.res(r12_88),.clk(clk),.wout(w12_88));
	PE pe12_89(.x(x89),.w(w12_88),.acc(r12_88),.res(r12_89),.clk(clk),.wout(w12_89));
	PE pe12_90(.x(x90),.w(w12_89),.acc(r12_89),.res(r12_90),.clk(clk),.wout(w12_90));
	PE pe12_91(.x(x91),.w(w12_90),.acc(r12_90),.res(r12_91),.clk(clk),.wout(w12_91));
	PE pe12_92(.x(x92),.w(w12_91),.acc(r12_91),.res(r12_92),.clk(clk),.wout(w12_92));
	PE pe12_93(.x(x93),.w(w12_92),.acc(r12_92),.res(r12_93),.clk(clk),.wout(w12_93));
	PE pe12_94(.x(x94),.w(w12_93),.acc(r12_93),.res(r12_94),.clk(clk),.wout(w12_94));
	PE pe12_95(.x(x95),.w(w12_94),.acc(r12_94),.res(r12_95),.clk(clk),.wout(w12_95));
	PE pe12_96(.x(x96),.w(w12_95),.acc(r12_95),.res(r12_96),.clk(clk),.wout(w12_96));
	PE pe12_97(.x(x97),.w(w12_96),.acc(r12_96),.res(r12_97),.clk(clk),.wout(w12_97));
	PE pe12_98(.x(x98),.w(w12_97),.acc(r12_97),.res(r12_98),.clk(clk),.wout(w12_98));
	PE pe12_99(.x(x99),.w(w12_98),.acc(r12_98),.res(r12_99),.clk(clk),.wout(w12_99));
	PE pe12_100(.x(x100),.w(w12_99),.acc(r12_99),.res(r12_100),.clk(clk),.wout(w12_100));
	PE pe12_101(.x(x101),.w(w12_100),.acc(r12_100),.res(r12_101),.clk(clk),.wout(w12_101));
	PE pe12_102(.x(x102),.w(w12_101),.acc(r12_101),.res(r12_102),.clk(clk),.wout(w12_102));
	PE pe12_103(.x(x103),.w(w12_102),.acc(r12_102),.res(r12_103),.clk(clk),.wout(w12_103));
	PE pe12_104(.x(x104),.w(w12_103),.acc(r12_103),.res(r12_104),.clk(clk),.wout(w12_104));
	PE pe12_105(.x(x105),.w(w12_104),.acc(r12_104),.res(r12_105),.clk(clk),.wout(w12_105));
	PE pe12_106(.x(x106),.w(w12_105),.acc(r12_105),.res(r12_106),.clk(clk),.wout(w12_106));
	PE pe12_107(.x(x107),.w(w12_106),.acc(r12_106),.res(r12_107),.clk(clk),.wout(w12_107));
	PE pe12_108(.x(x108),.w(w12_107),.acc(r12_107),.res(r12_108),.clk(clk),.wout(w12_108));
	PE pe12_109(.x(x109),.w(w12_108),.acc(r12_108),.res(r12_109),.clk(clk),.wout(w12_109));
	PE pe12_110(.x(x110),.w(w12_109),.acc(r12_109),.res(r12_110),.clk(clk),.wout(w12_110));
	PE pe12_111(.x(x111),.w(w12_110),.acc(r12_110),.res(r12_111),.clk(clk),.wout(w12_111));
	PE pe12_112(.x(x112),.w(w12_111),.acc(r12_111),.res(r12_112),.clk(clk),.wout(w12_112));
	PE pe12_113(.x(x113),.w(w12_112),.acc(r12_112),.res(r12_113),.clk(clk),.wout(w12_113));
	PE pe12_114(.x(x114),.w(w12_113),.acc(r12_113),.res(r12_114),.clk(clk),.wout(w12_114));
	PE pe12_115(.x(x115),.w(w12_114),.acc(r12_114),.res(r12_115),.clk(clk),.wout(w12_115));
	PE pe12_116(.x(x116),.w(w12_115),.acc(r12_115),.res(r12_116),.clk(clk),.wout(w12_116));
	PE pe12_117(.x(x117),.w(w12_116),.acc(r12_116),.res(r12_117),.clk(clk),.wout(w12_117));
	PE pe12_118(.x(x118),.w(w12_117),.acc(r12_117),.res(r12_118),.clk(clk),.wout(w12_118));
	PE pe12_119(.x(x119),.w(w12_118),.acc(r12_118),.res(r12_119),.clk(clk),.wout(w12_119));
	PE pe12_120(.x(x120),.w(w12_119),.acc(r12_119),.res(r12_120),.clk(clk),.wout(w12_120));
	PE pe12_121(.x(x121),.w(w12_120),.acc(r12_120),.res(r12_121),.clk(clk),.wout(w12_121));
	PE pe12_122(.x(x122),.w(w12_121),.acc(r12_121),.res(r12_122),.clk(clk),.wout(w12_122));
	PE pe12_123(.x(x123),.w(w12_122),.acc(r12_122),.res(r12_123),.clk(clk),.wout(w12_123));
	PE pe12_124(.x(x124),.w(w12_123),.acc(r12_123),.res(r12_124),.clk(clk),.wout(w12_124));
	PE pe12_125(.x(x125),.w(w12_124),.acc(r12_124),.res(r12_125),.clk(clk),.wout(w12_125));
	PE pe12_126(.x(x126),.w(w12_125),.acc(r12_125),.res(r12_126),.clk(clk),.wout(w12_126));
	PE pe12_127(.x(x127),.w(w12_126),.acc(r12_126),.res(result12),.clk(clk),.wout(weight12));

	PE pe13_0(.x(x0),.w(w13),.acc(32'h0),.res(r13_0),.clk(clk),.wout(w13_0));
	PE pe13_1(.x(x1),.w(w13_0),.acc(r13_0),.res(r13_1),.clk(clk),.wout(w13_1));
	PE pe13_2(.x(x2),.w(w13_1),.acc(r13_1),.res(r13_2),.clk(clk),.wout(w13_2));
	PE pe13_3(.x(x3),.w(w13_2),.acc(r13_2),.res(r13_3),.clk(clk),.wout(w13_3));
	PE pe13_4(.x(x4),.w(w13_3),.acc(r13_3),.res(r13_4),.clk(clk),.wout(w13_4));
	PE pe13_5(.x(x5),.w(w13_4),.acc(r13_4),.res(r13_5),.clk(clk),.wout(w13_5));
	PE pe13_6(.x(x6),.w(w13_5),.acc(r13_5),.res(r13_6),.clk(clk),.wout(w13_6));
	PE pe13_7(.x(x7),.w(w13_6),.acc(r13_6),.res(r13_7),.clk(clk),.wout(w13_7));
	PE pe13_8(.x(x8),.w(w13_7),.acc(r13_7),.res(r13_8),.clk(clk),.wout(w13_8));
	PE pe13_9(.x(x9),.w(w13_8),.acc(r13_8),.res(r13_9),.clk(clk),.wout(w13_9));
	PE pe13_10(.x(x10),.w(w13_9),.acc(r13_9),.res(r13_10),.clk(clk),.wout(w13_10));
	PE pe13_11(.x(x11),.w(w13_10),.acc(r13_10),.res(r13_11),.clk(clk),.wout(w13_11));
	PE pe13_12(.x(x12),.w(w13_11),.acc(r13_11),.res(r13_12),.clk(clk),.wout(w13_12));
	PE pe13_13(.x(x13),.w(w13_12),.acc(r13_12),.res(r13_13),.clk(clk),.wout(w13_13));
	PE pe13_14(.x(x14),.w(w13_13),.acc(r13_13),.res(r13_14),.clk(clk),.wout(w13_14));
	PE pe13_15(.x(x15),.w(w13_14),.acc(r13_14),.res(r13_15),.clk(clk),.wout(w13_15));
	PE pe13_16(.x(x16),.w(w13_15),.acc(r13_15),.res(r13_16),.clk(clk),.wout(w13_16));
	PE pe13_17(.x(x17),.w(w13_16),.acc(r13_16),.res(r13_17),.clk(clk),.wout(w13_17));
	PE pe13_18(.x(x18),.w(w13_17),.acc(r13_17),.res(r13_18),.clk(clk),.wout(w13_18));
	PE pe13_19(.x(x19),.w(w13_18),.acc(r13_18),.res(r13_19),.clk(clk),.wout(w13_19));
	PE pe13_20(.x(x20),.w(w13_19),.acc(r13_19),.res(r13_20),.clk(clk),.wout(w13_20));
	PE pe13_21(.x(x21),.w(w13_20),.acc(r13_20),.res(r13_21),.clk(clk),.wout(w13_21));
	PE pe13_22(.x(x22),.w(w13_21),.acc(r13_21),.res(r13_22),.clk(clk),.wout(w13_22));
	PE pe13_23(.x(x23),.w(w13_22),.acc(r13_22),.res(r13_23),.clk(clk),.wout(w13_23));
	PE pe13_24(.x(x24),.w(w13_23),.acc(r13_23),.res(r13_24),.clk(clk),.wout(w13_24));
	PE pe13_25(.x(x25),.w(w13_24),.acc(r13_24),.res(r13_25),.clk(clk),.wout(w13_25));
	PE pe13_26(.x(x26),.w(w13_25),.acc(r13_25),.res(r13_26),.clk(clk),.wout(w13_26));
	PE pe13_27(.x(x27),.w(w13_26),.acc(r13_26),.res(r13_27),.clk(clk),.wout(w13_27));
	PE pe13_28(.x(x28),.w(w13_27),.acc(r13_27),.res(r13_28),.clk(clk),.wout(w13_28));
	PE pe13_29(.x(x29),.w(w13_28),.acc(r13_28),.res(r13_29),.clk(clk),.wout(w13_29));
	PE pe13_30(.x(x30),.w(w13_29),.acc(r13_29),.res(r13_30),.clk(clk),.wout(w13_30));
	PE pe13_31(.x(x31),.w(w13_30),.acc(r13_30),.res(r13_31),.clk(clk),.wout(w13_31));
	PE pe13_32(.x(x32),.w(w13_31),.acc(r13_31),.res(r13_32),.clk(clk),.wout(w13_32));
	PE pe13_33(.x(x33),.w(w13_32),.acc(r13_32),.res(r13_33),.clk(clk),.wout(w13_33));
	PE pe13_34(.x(x34),.w(w13_33),.acc(r13_33),.res(r13_34),.clk(clk),.wout(w13_34));
	PE pe13_35(.x(x35),.w(w13_34),.acc(r13_34),.res(r13_35),.clk(clk),.wout(w13_35));
	PE pe13_36(.x(x36),.w(w13_35),.acc(r13_35),.res(r13_36),.clk(clk),.wout(w13_36));
	PE pe13_37(.x(x37),.w(w13_36),.acc(r13_36),.res(r13_37),.clk(clk),.wout(w13_37));
	PE pe13_38(.x(x38),.w(w13_37),.acc(r13_37),.res(r13_38),.clk(clk),.wout(w13_38));
	PE pe13_39(.x(x39),.w(w13_38),.acc(r13_38),.res(r13_39),.clk(clk),.wout(w13_39));
	PE pe13_40(.x(x40),.w(w13_39),.acc(r13_39),.res(r13_40),.clk(clk),.wout(w13_40));
	PE pe13_41(.x(x41),.w(w13_40),.acc(r13_40),.res(r13_41),.clk(clk),.wout(w13_41));
	PE pe13_42(.x(x42),.w(w13_41),.acc(r13_41),.res(r13_42),.clk(clk),.wout(w13_42));
	PE pe13_43(.x(x43),.w(w13_42),.acc(r13_42),.res(r13_43),.clk(clk),.wout(w13_43));
	PE pe13_44(.x(x44),.w(w13_43),.acc(r13_43),.res(r13_44),.clk(clk),.wout(w13_44));
	PE pe13_45(.x(x45),.w(w13_44),.acc(r13_44),.res(r13_45),.clk(clk),.wout(w13_45));
	PE pe13_46(.x(x46),.w(w13_45),.acc(r13_45),.res(r13_46),.clk(clk),.wout(w13_46));
	PE pe13_47(.x(x47),.w(w13_46),.acc(r13_46),.res(r13_47),.clk(clk),.wout(w13_47));
	PE pe13_48(.x(x48),.w(w13_47),.acc(r13_47),.res(r13_48),.clk(clk),.wout(w13_48));
	PE pe13_49(.x(x49),.w(w13_48),.acc(r13_48),.res(r13_49),.clk(clk),.wout(w13_49));
	PE pe13_50(.x(x50),.w(w13_49),.acc(r13_49),.res(r13_50),.clk(clk),.wout(w13_50));
	PE pe13_51(.x(x51),.w(w13_50),.acc(r13_50),.res(r13_51),.clk(clk),.wout(w13_51));
	PE pe13_52(.x(x52),.w(w13_51),.acc(r13_51),.res(r13_52),.clk(clk),.wout(w13_52));
	PE pe13_53(.x(x53),.w(w13_52),.acc(r13_52),.res(r13_53),.clk(clk),.wout(w13_53));
	PE pe13_54(.x(x54),.w(w13_53),.acc(r13_53),.res(r13_54),.clk(clk),.wout(w13_54));
	PE pe13_55(.x(x55),.w(w13_54),.acc(r13_54),.res(r13_55),.clk(clk),.wout(w13_55));
	PE pe13_56(.x(x56),.w(w13_55),.acc(r13_55),.res(r13_56),.clk(clk),.wout(w13_56));
	PE pe13_57(.x(x57),.w(w13_56),.acc(r13_56),.res(r13_57),.clk(clk),.wout(w13_57));
	PE pe13_58(.x(x58),.w(w13_57),.acc(r13_57),.res(r13_58),.clk(clk),.wout(w13_58));
	PE pe13_59(.x(x59),.w(w13_58),.acc(r13_58),.res(r13_59),.clk(clk),.wout(w13_59));
	PE pe13_60(.x(x60),.w(w13_59),.acc(r13_59),.res(r13_60),.clk(clk),.wout(w13_60));
	PE pe13_61(.x(x61),.w(w13_60),.acc(r13_60),.res(r13_61),.clk(clk),.wout(w13_61));
	PE pe13_62(.x(x62),.w(w13_61),.acc(r13_61),.res(r13_62),.clk(clk),.wout(w13_62));
	PE pe13_63(.x(x63),.w(w13_62),.acc(r13_62),.res(r13_63),.clk(clk),.wout(w13_63));
	PE pe13_64(.x(x64),.w(w13_63),.acc(r13_63),.res(r13_64),.clk(clk),.wout(w13_64));
	PE pe13_65(.x(x65),.w(w13_64),.acc(r13_64),.res(r13_65),.clk(clk),.wout(w13_65));
	PE pe13_66(.x(x66),.w(w13_65),.acc(r13_65),.res(r13_66),.clk(clk),.wout(w13_66));
	PE pe13_67(.x(x67),.w(w13_66),.acc(r13_66),.res(r13_67),.clk(clk),.wout(w13_67));
	PE pe13_68(.x(x68),.w(w13_67),.acc(r13_67),.res(r13_68),.clk(clk),.wout(w13_68));
	PE pe13_69(.x(x69),.w(w13_68),.acc(r13_68),.res(r13_69),.clk(clk),.wout(w13_69));
	PE pe13_70(.x(x70),.w(w13_69),.acc(r13_69),.res(r13_70),.clk(clk),.wout(w13_70));
	PE pe13_71(.x(x71),.w(w13_70),.acc(r13_70),.res(r13_71),.clk(clk),.wout(w13_71));
	PE pe13_72(.x(x72),.w(w13_71),.acc(r13_71),.res(r13_72),.clk(clk),.wout(w13_72));
	PE pe13_73(.x(x73),.w(w13_72),.acc(r13_72),.res(r13_73),.clk(clk),.wout(w13_73));
	PE pe13_74(.x(x74),.w(w13_73),.acc(r13_73),.res(r13_74),.clk(clk),.wout(w13_74));
	PE pe13_75(.x(x75),.w(w13_74),.acc(r13_74),.res(r13_75),.clk(clk),.wout(w13_75));
	PE pe13_76(.x(x76),.w(w13_75),.acc(r13_75),.res(r13_76),.clk(clk),.wout(w13_76));
	PE pe13_77(.x(x77),.w(w13_76),.acc(r13_76),.res(r13_77),.clk(clk),.wout(w13_77));
	PE pe13_78(.x(x78),.w(w13_77),.acc(r13_77),.res(r13_78),.clk(clk),.wout(w13_78));
	PE pe13_79(.x(x79),.w(w13_78),.acc(r13_78),.res(r13_79),.clk(clk),.wout(w13_79));
	PE pe13_80(.x(x80),.w(w13_79),.acc(r13_79),.res(r13_80),.clk(clk),.wout(w13_80));
	PE pe13_81(.x(x81),.w(w13_80),.acc(r13_80),.res(r13_81),.clk(clk),.wout(w13_81));
	PE pe13_82(.x(x82),.w(w13_81),.acc(r13_81),.res(r13_82),.clk(clk),.wout(w13_82));
	PE pe13_83(.x(x83),.w(w13_82),.acc(r13_82),.res(r13_83),.clk(clk),.wout(w13_83));
	PE pe13_84(.x(x84),.w(w13_83),.acc(r13_83),.res(r13_84),.clk(clk),.wout(w13_84));
	PE pe13_85(.x(x85),.w(w13_84),.acc(r13_84),.res(r13_85),.clk(clk),.wout(w13_85));
	PE pe13_86(.x(x86),.w(w13_85),.acc(r13_85),.res(r13_86),.clk(clk),.wout(w13_86));
	PE pe13_87(.x(x87),.w(w13_86),.acc(r13_86),.res(r13_87),.clk(clk),.wout(w13_87));
	PE pe13_88(.x(x88),.w(w13_87),.acc(r13_87),.res(r13_88),.clk(clk),.wout(w13_88));
	PE pe13_89(.x(x89),.w(w13_88),.acc(r13_88),.res(r13_89),.clk(clk),.wout(w13_89));
	PE pe13_90(.x(x90),.w(w13_89),.acc(r13_89),.res(r13_90),.clk(clk),.wout(w13_90));
	PE pe13_91(.x(x91),.w(w13_90),.acc(r13_90),.res(r13_91),.clk(clk),.wout(w13_91));
	PE pe13_92(.x(x92),.w(w13_91),.acc(r13_91),.res(r13_92),.clk(clk),.wout(w13_92));
	PE pe13_93(.x(x93),.w(w13_92),.acc(r13_92),.res(r13_93),.clk(clk),.wout(w13_93));
	PE pe13_94(.x(x94),.w(w13_93),.acc(r13_93),.res(r13_94),.clk(clk),.wout(w13_94));
	PE pe13_95(.x(x95),.w(w13_94),.acc(r13_94),.res(r13_95),.clk(clk),.wout(w13_95));
	PE pe13_96(.x(x96),.w(w13_95),.acc(r13_95),.res(r13_96),.clk(clk),.wout(w13_96));
	PE pe13_97(.x(x97),.w(w13_96),.acc(r13_96),.res(r13_97),.clk(clk),.wout(w13_97));
	PE pe13_98(.x(x98),.w(w13_97),.acc(r13_97),.res(r13_98),.clk(clk),.wout(w13_98));
	PE pe13_99(.x(x99),.w(w13_98),.acc(r13_98),.res(r13_99),.clk(clk),.wout(w13_99));
	PE pe13_100(.x(x100),.w(w13_99),.acc(r13_99),.res(r13_100),.clk(clk),.wout(w13_100));
	PE pe13_101(.x(x101),.w(w13_100),.acc(r13_100),.res(r13_101),.clk(clk),.wout(w13_101));
	PE pe13_102(.x(x102),.w(w13_101),.acc(r13_101),.res(r13_102),.clk(clk),.wout(w13_102));
	PE pe13_103(.x(x103),.w(w13_102),.acc(r13_102),.res(r13_103),.clk(clk),.wout(w13_103));
	PE pe13_104(.x(x104),.w(w13_103),.acc(r13_103),.res(r13_104),.clk(clk),.wout(w13_104));
	PE pe13_105(.x(x105),.w(w13_104),.acc(r13_104),.res(r13_105),.clk(clk),.wout(w13_105));
	PE pe13_106(.x(x106),.w(w13_105),.acc(r13_105),.res(r13_106),.clk(clk),.wout(w13_106));
	PE pe13_107(.x(x107),.w(w13_106),.acc(r13_106),.res(r13_107),.clk(clk),.wout(w13_107));
	PE pe13_108(.x(x108),.w(w13_107),.acc(r13_107),.res(r13_108),.clk(clk),.wout(w13_108));
	PE pe13_109(.x(x109),.w(w13_108),.acc(r13_108),.res(r13_109),.clk(clk),.wout(w13_109));
	PE pe13_110(.x(x110),.w(w13_109),.acc(r13_109),.res(r13_110),.clk(clk),.wout(w13_110));
	PE pe13_111(.x(x111),.w(w13_110),.acc(r13_110),.res(r13_111),.clk(clk),.wout(w13_111));
	PE pe13_112(.x(x112),.w(w13_111),.acc(r13_111),.res(r13_112),.clk(clk),.wout(w13_112));
	PE pe13_113(.x(x113),.w(w13_112),.acc(r13_112),.res(r13_113),.clk(clk),.wout(w13_113));
	PE pe13_114(.x(x114),.w(w13_113),.acc(r13_113),.res(r13_114),.clk(clk),.wout(w13_114));
	PE pe13_115(.x(x115),.w(w13_114),.acc(r13_114),.res(r13_115),.clk(clk),.wout(w13_115));
	PE pe13_116(.x(x116),.w(w13_115),.acc(r13_115),.res(r13_116),.clk(clk),.wout(w13_116));
	PE pe13_117(.x(x117),.w(w13_116),.acc(r13_116),.res(r13_117),.clk(clk),.wout(w13_117));
	PE pe13_118(.x(x118),.w(w13_117),.acc(r13_117),.res(r13_118),.clk(clk),.wout(w13_118));
	PE pe13_119(.x(x119),.w(w13_118),.acc(r13_118),.res(r13_119),.clk(clk),.wout(w13_119));
	PE pe13_120(.x(x120),.w(w13_119),.acc(r13_119),.res(r13_120),.clk(clk),.wout(w13_120));
	PE pe13_121(.x(x121),.w(w13_120),.acc(r13_120),.res(r13_121),.clk(clk),.wout(w13_121));
	PE pe13_122(.x(x122),.w(w13_121),.acc(r13_121),.res(r13_122),.clk(clk),.wout(w13_122));
	PE pe13_123(.x(x123),.w(w13_122),.acc(r13_122),.res(r13_123),.clk(clk),.wout(w13_123));
	PE pe13_124(.x(x124),.w(w13_123),.acc(r13_123),.res(r13_124),.clk(clk),.wout(w13_124));
	PE pe13_125(.x(x125),.w(w13_124),.acc(r13_124),.res(r13_125),.clk(clk),.wout(w13_125));
	PE pe13_126(.x(x126),.w(w13_125),.acc(r13_125),.res(r13_126),.clk(clk),.wout(w13_126));
	PE pe13_127(.x(x127),.w(w13_126),.acc(r13_126),.res(result13),.clk(clk),.wout(weight13));

	PE pe14_0(.x(x0),.w(w14),.acc(32'h0),.res(r14_0),.clk(clk),.wout(w14_0));
	PE pe14_1(.x(x1),.w(w14_0),.acc(r14_0),.res(r14_1),.clk(clk),.wout(w14_1));
	PE pe14_2(.x(x2),.w(w14_1),.acc(r14_1),.res(r14_2),.clk(clk),.wout(w14_2));
	PE pe14_3(.x(x3),.w(w14_2),.acc(r14_2),.res(r14_3),.clk(clk),.wout(w14_3));
	PE pe14_4(.x(x4),.w(w14_3),.acc(r14_3),.res(r14_4),.clk(clk),.wout(w14_4));
	PE pe14_5(.x(x5),.w(w14_4),.acc(r14_4),.res(r14_5),.clk(clk),.wout(w14_5));
	PE pe14_6(.x(x6),.w(w14_5),.acc(r14_5),.res(r14_6),.clk(clk),.wout(w14_6));
	PE pe14_7(.x(x7),.w(w14_6),.acc(r14_6),.res(r14_7),.clk(clk),.wout(w14_7));
	PE pe14_8(.x(x8),.w(w14_7),.acc(r14_7),.res(r14_8),.clk(clk),.wout(w14_8));
	PE pe14_9(.x(x9),.w(w14_8),.acc(r14_8),.res(r14_9),.clk(clk),.wout(w14_9));
	PE pe14_10(.x(x10),.w(w14_9),.acc(r14_9),.res(r14_10),.clk(clk),.wout(w14_10));
	PE pe14_11(.x(x11),.w(w14_10),.acc(r14_10),.res(r14_11),.clk(clk),.wout(w14_11));
	PE pe14_12(.x(x12),.w(w14_11),.acc(r14_11),.res(r14_12),.clk(clk),.wout(w14_12));
	PE pe14_13(.x(x13),.w(w14_12),.acc(r14_12),.res(r14_13),.clk(clk),.wout(w14_13));
	PE pe14_14(.x(x14),.w(w14_13),.acc(r14_13),.res(r14_14),.clk(clk),.wout(w14_14));
	PE pe14_15(.x(x15),.w(w14_14),.acc(r14_14),.res(r14_15),.clk(clk),.wout(w14_15));
	PE pe14_16(.x(x16),.w(w14_15),.acc(r14_15),.res(r14_16),.clk(clk),.wout(w14_16));
	PE pe14_17(.x(x17),.w(w14_16),.acc(r14_16),.res(r14_17),.clk(clk),.wout(w14_17));
	PE pe14_18(.x(x18),.w(w14_17),.acc(r14_17),.res(r14_18),.clk(clk),.wout(w14_18));
	PE pe14_19(.x(x19),.w(w14_18),.acc(r14_18),.res(r14_19),.clk(clk),.wout(w14_19));
	PE pe14_20(.x(x20),.w(w14_19),.acc(r14_19),.res(r14_20),.clk(clk),.wout(w14_20));
	PE pe14_21(.x(x21),.w(w14_20),.acc(r14_20),.res(r14_21),.clk(clk),.wout(w14_21));
	PE pe14_22(.x(x22),.w(w14_21),.acc(r14_21),.res(r14_22),.clk(clk),.wout(w14_22));
	PE pe14_23(.x(x23),.w(w14_22),.acc(r14_22),.res(r14_23),.clk(clk),.wout(w14_23));
	PE pe14_24(.x(x24),.w(w14_23),.acc(r14_23),.res(r14_24),.clk(clk),.wout(w14_24));
	PE pe14_25(.x(x25),.w(w14_24),.acc(r14_24),.res(r14_25),.clk(clk),.wout(w14_25));
	PE pe14_26(.x(x26),.w(w14_25),.acc(r14_25),.res(r14_26),.clk(clk),.wout(w14_26));
	PE pe14_27(.x(x27),.w(w14_26),.acc(r14_26),.res(r14_27),.clk(clk),.wout(w14_27));
	PE pe14_28(.x(x28),.w(w14_27),.acc(r14_27),.res(r14_28),.clk(clk),.wout(w14_28));
	PE pe14_29(.x(x29),.w(w14_28),.acc(r14_28),.res(r14_29),.clk(clk),.wout(w14_29));
	PE pe14_30(.x(x30),.w(w14_29),.acc(r14_29),.res(r14_30),.clk(clk),.wout(w14_30));
	PE pe14_31(.x(x31),.w(w14_30),.acc(r14_30),.res(r14_31),.clk(clk),.wout(w14_31));
	PE pe14_32(.x(x32),.w(w14_31),.acc(r14_31),.res(r14_32),.clk(clk),.wout(w14_32));
	PE pe14_33(.x(x33),.w(w14_32),.acc(r14_32),.res(r14_33),.clk(clk),.wout(w14_33));
	PE pe14_34(.x(x34),.w(w14_33),.acc(r14_33),.res(r14_34),.clk(clk),.wout(w14_34));
	PE pe14_35(.x(x35),.w(w14_34),.acc(r14_34),.res(r14_35),.clk(clk),.wout(w14_35));
	PE pe14_36(.x(x36),.w(w14_35),.acc(r14_35),.res(r14_36),.clk(clk),.wout(w14_36));
	PE pe14_37(.x(x37),.w(w14_36),.acc(r14_36),.res(r14_37),.clk(clk),.wout(w14_37));
	PE pe14_38(.x(x38),.w(w14_37),.acc(r14_37),.res(r14_38),.clk(clk),.wout(w14_38));
	PE pe14_39(.x(x39),.w(w14_38),.acc(r14_38),.res(r14_39),.clk(clk),.wout(w14_39));
	PE pe14_40(.x(x40),.w(w14_39),.acc(r14_39),.res(r14_40),.clk(clk),.wout(w14_40));
	PE pe14_41(.x(x41),.w(w14_40),.acc(r14_40),.res(r14_41),.clk(clk),.wout(w14_41));
	PE pe14_42(.x(x42),.w(w14_41),.acc(r14_41),.res(r14_42),.clk(clk),.wout(w14_42));
	PE pe14_43(.x(x43),.w(w14_42),.acc(r14_42),.res(r14_43),.clk(clk),.wout(w14_43));
	PE pe14_44(.x(x44),.w(w14_43),.acc(r14_43),.res(r14_44),.clk(clk),.wout(w14_44));
	PE pe14_45(.x(x45),.w(w14_44),.acc(r14_44),.res(r14_45),.clk(clk),.wout(w14_45));
	PE pe14_46(.x(x46),.w(w14_45),.acc(r14_45),.res(r14_46),.clk(clk),.wout(w14_46));
	PE pe14_47(.x(x47),.w(w14_46),.acc(r14_46),.res(r14_47),.clk(clk),.wout(w14_47));
	PE pe14_48(.x(x48),.w(w14_47),.acc(r14_47),.res(r14_48),.clk(clk),.wout(w14_48));
	PE pe14_49(.x(x49),.w(w14_48),.acc(r14_48),.res(r14_49),.clk(clk),.wout(w14_49));
	PE pe14_50(.x(x50),.w(w14_49),.acc(r14_49),.res(r14_50),.clk(clk),.wout(w14_50));
	PE pe14_51(.x(x51),.w(w14_50),.acc(r14_50),.res(r14_51),.clk(clk),.wout(w14_51));
	PE pe14_52(.x(x52),.w(w14_51),.acc(r14_51),.res(r14_52),.clk(clk),.wout(w14_52));
	PE pe14_53(.x(x53),.w(w14_52),.acc(r14_52),.res(r14_53),.clk(clk),.wout(w14_53));
	PE pe14_54(.x(x54),.w(w14_53),.acc(r14_53),.res(r14_54),.clk(clk),.wout(w14_54));
	PE pe14_55(.x(x55),.w(w14_54),.acc(r14_54),.res(r14_55),.clk(clk),.wout(w14_55));
	PE pe14_56(.x(x56),.w(w14_55),.acc(r14_55),.res(r14_56),.clk(clk),.wout(w14_56));
	PE pe14_57(.x(x57),.w(w14_56),.acc(r14_56),.res(r14_57),.clk(clk),.wout(w14_57));
	PE pe14_58(.x(x58),.w(w14_57),.acc(r14_57),.res(r14_58),.clk(clk),.wout(w14_58));
	PE pe14_59(.x(x59),.w(w14_58),.acc(r14_58),.res(r14_59),.clk(clk),.wout(w14_59));
	PE pe14_60(.x(x60),.w(w14_59),.acc(r14_59),.res(r14_60),.clk(clk),.wout(w14_60));
	PE pe14_61(.x(x61),.w(w14_60),.acc(r14_60),.res(r14_61),.clk(clk),.wout(w14_61));
	PE pe14_62(.x(x62),.w(w14_61),.acc(r14_61),.res(r14_62),.clk(clk),.wout(w14_62));
	PE pe14_63(.x(x63),.w(w14_62),.acc(r14_62),.res(r14_63),.clk(clk),.wout(w14_63));
	PE pe14_64(.x(x64),.w(w14_63),.acc(r14_63),.res(r14_64),.clk(clk),.wout(w14_64));
	PE pe14_65(.x(x65),.w(w14_64),.acc(r14_64),.res(r14_65),.clk(clk),.wout(w14_65));
	PE pe14_66(.x(x66),.w(w14_65),.acc(r14_65),.res(r14_66),.clk(clk),.wout(w14_66));
	PE pe14_67(.x(x67),.w(w14_66),.acc(r14_66),.res(r14_67),.clk(clk),.wout(w14_67));
	PE pe14_68(.x(x68),.w(w14_67),.acc(r14_67),.res(r14_68),.clk(clk),.wout(w14_68));
	PE pe14_69(.x(x69),.w(w14_68),.acc(r14_68),.res(r14_69),.clk(clk),.wout(w14_69));
	PE pe14_70(.x(x70),.w(w14_69),.acc(r14_69),.res(r14_70),.clk(clk),.wout(w14_70));
	PE pe14_71(.x(x71),.w(w14_70),.acc(r14_70),.res(r14_71),.clk(clk),.wout(w14_71));
	PE pe14_72(.x(x72),.w(w14_71),.acc(r14_71),.res(r14_72),.clk(clk),.wout(w14_72));
	PE pe14_73(.x(x73),.w(w14_72),.acc(r14_72),.res(r14_73),.clk(clk),.wout(w14_73));
	PE pe14_74(.x(x74),.w(w14_73),.acc(r14_73),.res(r14_74),.clk(clk),.wout(w14_74));
	PE pe14_75(.x(x75),.w(w14_74),.acc(r14_74),.res(r14_75),.clk(clk),.wout(w14_75));
	PE pe14_76(.x(x76),.w(w14_75),.acc(r14_75),.res(r14_76),.clk(clk),.wout(w14_76));
	PE pe14_77(.x(x77),.w(w14_76),.acc(r14_76),.res(r14_77),.clk(clk),.wout(w14_77));
	PE pe14_78(.x(x78),.w(w14_77),.acc(r14_77),.res(r14_78),.clk(clk),.wout(w14_78));
	PE pe14_79(.x(x79),.w(w14_78),.acc(r14_78),.res(r14_79),.clk(clk),.wout(w14_79));
	PE pe14_80(.x(x80),.w(w14_79),.acc(r14_79),.res(r14_80),.clk(clk),.wout(w14_80));
	PE pe14_81(.x(x81),.w(w14_80),.acc(r14_80),.res(r14_81),.clk(clk),.wout(w14_81));
	PE pe14_82(.x(x82),.w(w14_81),.acc(r14_81),.res(r14_82),.clk(clk),.wout(w14_82));
	PE pe14_83(.x(x83),.w(w14_82),.acc(r14_82),.res(r14_83),.clk(clk),.wout(w14_83));
	PE pe14_84(.x(x84),.w(w14_83),.acc(r14_83),.res(r14_84),.clk(clk),.wout(w14_84));
	PE pe14_85(.x(x85),.w(w14_84),.acc(r14_84),.res(r14_85),.clk(clk),.wout(w14_85));
	PE pe14_86(.x(x86),.w(w14_85),.acc(r14_85),.res(r14_86),.clk(clk),.wout(w14_86));
	PE pe14_87(.x(x87),.w(w14_86),.acc(r14_86),.res(r14_87),.clk(clk),.wout(w14_87));
	PE pe14_88(.x(x88),.w(w14_87),.acc(r14_87),.res(r14_88),.clk(clk),.wout(w14_88));
	PE pe14_89(.x(x89),.w(w14_88),.acc(r14_88),.res(r14_89),.clk(clk),.wout(w14_89));
	PE pe14_90(.x(x90),.w(w14_89),.acc(r14_89),.res(r14_90),.clk(clk),.wout(w14_90));
	PE pe14_91(.x(x91),.w(w14_90),.acc(r14_90),.res(r14_91),.clk(clk),.wout(w14_91));
	PE pe14_92(.x(x92),.w(w14_91),.acc(r14_91),.res(r14_92),.clk(clk),.wout(w14_92));
	PE pe14_93(.x(x93),.w(w14_92),.acc(r14_92),.res(r14_93),.clk(clk),.wout(w14_93));
	PE pe14_94(.x(x94),.w(w14_93),.acc(r14_93),.res(r14_94),.clk(clk),.wout(w14_94));
	PE pe14_95(.x(x95),.w(w14_94),.acc(r14_94),.res(r14_95),.clk(clk),.wout(w14_95));
	PE pe14_96(.x(x96),.w(w14_95),.acc(r14_95),.res(r14_96),.clk(clk),.wout(w14_96));
	PE pe14_97(.x(x97),.w(w14_96),.acc(r14_96),.res(r14_97),.clk(clk),.wout(w14_97));
	PE pe14_98(.x(x98),.w(w14_97),.acc(r14_97),.res(r14_98),.clk(clk),.wout(w14_98));
	PE pe14_99(.x(x99),.w(w14_98),.acc(r14_98),.res(r14_99),.clk(clk),.wout(w14_99));
	PE pe14_100(.x(x100),.w(w14_99),.acc(r14_99),.res(r14_100),.clk(clk),.wout(w14_100));
	PE pe14_101(.x(x101),.w(w14_100),.acc(r14_100),.res(r14_101),.clk(clk),.wout(w14_101));
	PE pe14_102(.x(x102),.w(w14_101),.acc(r14_101),.res(r14_102),.clk(clk),.wout(w14_102));
	PE pe14_103(.x(x103),.w(w14_102),.acc(r14_102),.res(r14_103),.clk(clk),.wout(w14_103));
	PE pe14_104(.x(x104),.w(w14_103),.acc(r14_103),.res(r14_104),.clk(clk),.wout(w14_104));
	PE pe14_105(.x(x105),.w(w14_104),.acc(r14_104),.res(r14_105),.clk(clk),.wout(w14_105));
	PE pe14_106(.x(x106),.w(w14_105),.acc(r14_105),.res(r14_106),.clk(clk),.wout(w14_106));
	PE pe14_107(.x(x107),.w(w14_106),.acc(r14_106),.res(r14_107),.clk(clk),.wout(w14_107));
	PE pe14_108(.x(x108),.w(w14_107),.acc(r14_107),.res(r14_108),.clk(clk),.wout(w14_108));
	PE pe14_109(.x(x109),.w(w14_108),.acc(r14_108),.res(r14_109),.clk(clk),.wout(w14_109));
	PE pe14_110(.x(x110),.w(w14_109),.acc(r14_109),.res(r14_110),.clk(clk),.wout(w14_110));
	PE pe14_111(.x(x111),.w(w14_110),.acc(r14_110),.res(r14_111),.clk(clk),.wout(w14_111));
	PE pe14_112(.x(x112),.w(w14_111),.acc(r14_111),.res(r14_112),.clk(clk),.wout(w14_112));
	PE pe14_113(.x(x113),.w(w14_112),.acc(r14_112),.res(r14_113),.clk(clk),.wout(w14_113));
	PE pe14_114(.x(x114),.w(w14_113),.acc(r14_113),.res(r14_114),.clk(clk),.wout(w14_114));
	PE pe14_115(.x(x115),.w(w14_114),.acc(r14_114),.res(r14_115),.clk(clk),.wout(w14_115));
	PE pe14_116(.x(x116),.w(w14_115),.acc(r14_115),.res(r14_116),.clk(clk),.wout(w14_116));
	PE pe14_117(.x(x117),.w(w14_116),.acc(r14_116),.res(r14_117),.clk(clk),.wout(w14_117));
	PE pe14_118(.x(x118),.w(w14_117),.acc(r14_117),.res(r14_118),.clk(clk),.wout(w14_118));
	PE pe14_119(.x(x119),.w(w14_118),.acc(r14_118),.res(r14_119),.clk(clk),.wout(w14_119));
	PE pe14_120(.x(x120),.w(w14_119),.acc(r14_119),.res(r14_120),.clk(clk),.wout(w14_120));
	PE pe14_121(.x(x121),.w(w14_120),.acc(r14_120),.res(r14_121),.clk(clk),.wout(w14_121));
	PE pe14_122(.x(x122),.w(w14_121),.acc(r14_121),.res(r14_122),.clk(clk),.wout(w14_122));
	PE pe14_123(.x(x123),.w(w14_122),.acc(r14_122),.res(r14_123),.clk(clk),.wout(w14_123));
	PE pe14_124(.x(x124),.w(w14_123),.acc(r14_123),.res(r14_124),.clk(clk),.wout(w14_124));
	PE pe14_125(.x(x125),.w(w14_124),.acc(r14_124),.res(r14_125),.clk(clk),.wout(w14_125));
	PE pe14_126(.x(x126),.w(w14_125),.acc(r14_125),.res(r14_126),.clk(clk),.wout(w14_126));
	PE pe14_127(.x(x127),.w(w14_126),.acc(r14_126),.res(result14),.clk(clk),.wout(weight14));

	PE pe15_0(.x(x0),.w(w15),.acc(32'h0),.res(r15_0),.clk(clk),.wout(w15_0));
	PE pe15_1(.x(x1),.w(w15_0),.acc(r15_0),.res(r15_1),.clk(clk),.wout(w15_1));
	PE pe15_2(.x(x2),.w(w15_1),.acc(r15_1),.res(r15_2),.clk(clk),.wout(w15_2));
	PE pe15_3(.x(x3),.w(w15_2),.acc(r15_2),.res(r15_3),.clk(clk),.wout(w15_3));
	PE pe15_4(.x(x4),.w(w15_3),.acc(r15_3),.res(r15_4),.clk(clk),.wout(w15_4));
	PE pe15_5(.x(x5),.w(w15_4),.acc(r15_4),.res(r15_5),.clk(clk),.wout(w15_5));
	PE pe15_6(.x(x6),.w(w15_5),.acc(r15_5),.res(r15_6),.clk(clk),.wout(w15_6));
	PE pe15_7(.x(x7),.w(w15_6),.acc(r15_6),.res(r15_7),.clk(clk),.wout(w15_7));
	PE pe15_8(.x(x8),.w(w15_7),.acc(r15_7),.res(r15_8),.clk(clk),.wout(w15_8));
	PE pe15_9(.x(x9),.w(w15_8),.acc(r15_8),.res(r15_9),.clk(clk),.wout(w15_9));
	PE pe15_10(.x(x10),.w(w15_9),.acc(r15_9),.res(r15_10),.clk(clk),.wout(w15_10));
	PE pe15_11(.x(x11),.w(w15_10),.acc(r15_10),.res(r15_11),.clk(clk),.wout(w15_11));
	PE pe15_12(.x(x12),.w(w15_11),.acc(r15_11),.res(r15_12),.clk(clk),.wout(w15_12));
	PE pe15_13(.x(x13),.w(w15_12),.acc(r15_12),.res(r15_13),.clk(clk),.wout(w15_13));
	PE pe15_14(.x(x14),.w(w15_13),.acc(r15_13),.res(r15_14),.clk(clk),.wout(w15_14));
	PE pe15_15(.x(x15),.w(w15_14),.acc(r15_14),.res(r15_15),.clk(clk),.wout(w15_15));
	PE pe15_16(.x(x16),.w(w15_15),.acc(r15_15),.res(r15_16),.clk(clk),.wout(w15_16));
	PE pe15_17(.x(x17),.w(w15_16),.acc(r15_16),.res(r15_17),.clk(clk),.wout(w15_17));
	PE pe15_18(.x(x18),.w(w15_17),.acc(r15_17),.res(r15_18),.clk(clk),.wout(w15_18));
	PE pe15_19(.x(x19),.w(w15_18),.acc(r15_18),.res(r15_19),.clk(clk),.wout(w15_19));
	PE pe15_20(.x(x20),.w(w15_19),.acc(r15_19),.res(r15_20),.clk(clk),.wout(w15_20));
	PE pe15_21(.x(x21),.w(w15_20),.acc(r15_20),.res(r15_21),.clk(clk),.wout(w15_21));
	PE pe15_22(.x(x22),.w(w15_21),.acc(r15_21),.res(r15_22),.clk(clk),.wout(w15_22));
	PE pe15_23(.x(x23),.w(w15_22),.acc(r15_22),.res(r15_23),.clk(clk),.wout(w15_23));
	PE pe15_24(.x(x24),.w(w15_23),.acc(r15_23),.res(r15_24),.clk(clk),.wout(w15_24));
	PE pe15_25(.x(x25),.w(w15_24),.acc(r15_24),.res(r15_25),.clk(clk),.wout(w15_25));
	PE pe15_26(.x(x26),.w(w15_25),.acc(r15_25),.res(r15_26),.clk(clk),.wout(w15_26));
	PE pe15_27(.x(x27),.w(w15_26),.acc(r15_26),.res(r15_27),.clk(clk),.wout(w15_27));
	PE pe15_28(.x(x28),.w(w15_27),.acc(r15_27),.res(r15_28),.clk(clk),.wout(w15_28));
	PE pe15_29(.x(x29),.w(w15_28),.acc(r15_28),.res(r15_29),.clk(clk),.wout(w15_29));
	PE pe15_30(.x(x30),.w(w15_29),.acc(r15_29),.res(r15_30),.clk(clk),.wout(w15_30));
	PE pe15_31(.x(x31),.w(w15_30),.acc(r15_30),.res(r15_31),.clk(clk),.wout(w15_31));
	PE pe15_32(.x(x32),.w(w15_31),.acc(r15_31),.res(r15_32),.clk(clk),.wout(w15_32));
	PE pe15_33(.x(x33),.w(w15_32),.acc(r15_32),.res(r15_33),.clk(clk),.wout(w15_33));
	PE pe15_34(.x(x34),.w(w15_33),.acc(r15_33),.res(r15_34),.clk(clk),.wout(w15_34));
	PE pe15_35(.x(x35),.w(w15_34),.acc(r15_34),.res(r15_35),.clk(clk),.wout(w15_35));
	PE pe15_36(.x(x36),.w(w15_35),.acc(r15_35),.res(r15_36),.clk(clk),.wout(w15_36));
	PE pe15_37(.x(x37),.w(w15_36),.acc(r15_36),.res(r15_37),.clk(clk),.wout(w15_37));
	PE pe15_38(.x(x38),.w(w15_37),.acc(r15_37),.res(r15_38),.clk(clk),.wout(w15_38));
	PE pe15_39(.x(x39),.w(w15_38),.acc(r15_38),.res(r15_39),.clk(clk),.wout(w15_39));
	PE pe15_40(.x(x40),.w(w15_39),.acc(r15_39),.res(r15_40),.clk(clk),.wout(w15_40));
	PE pe15_41(.x(x41),.w(w15_40),.acc(r15_40),.res(r15_41),.clk(clk),.wout(w15_41));
	PE pe15_42(.x(x42),.w(w15_41),.acc(r15_41),.res(r15_42),.clk(clk),.wout(w15_42));
	PE pe15_43(.x(x43),.w(w15_42),.acc(r15_42),.res(r15_43),.clk(clk),.wout(w15_43));
	PE pe15_44(.x(x44),.w(w15_43),.acc(r15_43),.res(r15_44),.clk(clk),.wout(w15_44));
	PE pe15_45(.x(x45),.w(w15_44),.acc(r15_44),.res(r15_45),.clk(clk),.wout(w15_45));
	PE pe15_46(.x(x46),.w(w15_45),.acc(r15_45),.res(r15_46),.clk(clk),.wout(w15_46));
	PE pe15_47(.x(x47),.w(w15_46),.acc(r15_46),.res(r15_47),.clk(clk),.wout(w15_47));
	PE pe15_48(.x(x48),.w(w15_47),.acc(r15_47),.res(r15_48),.clk(clk),.wout(w15_48));
	PE pe15_49(.x(x49),.w(w15_48),.acc(r15_48),.res(r15_49),.clk(clk),.wout(w15_49));
	PE pe15_50(.x(x50),.w(w15_49),.acc(r15_49),.res(r15_50),.clk(clk),.wout(w15_50));
	PE pe15_51(.x(x51),.w(w15_50),.acc(r15_50),.res(r15_51),.clk(clk),.wout(w15_51));
	PE pe15_52(.x(x52),.w(w15_51),.acc(r15_51),.res(r15_52),.clk(clk),.wout(w15_52));
	PE pe15_53(.x(x53),.w(w15_52),.acc(r15_52),.res(r15_53),.clk(clk),.wout(w15_53));
	PE pe15_54(.x(x54),.w(w15_53),.acc(r15_53),.res(r15_54),.clk(clk),.wout(w15_54));
	PE pe15_55(.x(x55),.w(w15_54),.acc(r15_54),.res(r15_55),.clk(clk),.wout(w15_55));
	PE pe15_56(.x(x56),.w(w15_55),.acc(r15_55),.res(r15_56),.clk(clk),.wout(w15_56));
	PE pe15_57(.x(x57),.w(w15_56),.acc(r15_56),.res(r15_57),.clk(clk),.wout(w15_57));
	PE pe15_58(.x(x58),.w(w15_57),.acc(r15_57),.res(r15_58),.clk(clk),.wout(w15_58));
	PE pe15_59(.x(x59),.w(w15_58),.acc(r15_58),.res(r15_59),.clk(clk),.wout(w15_59));
	PE pe15_60(.x(x60),.w(w15_59),.acc(r15_59),.res(r15_60),.clk(clk),.wout(w15_60));
	PE pe15_61(.x(x61),.w(w15_60),.acc(r15_60),.res(r15_61),.clk(clk),.wout(w15_61));
	PE pe15_62(.x(x62),.w(w15_61),.acc(r15_61),.res(r15_62),.clk(clk),.wout(w15_62));
	PE pe15_63(.x(x63),.w(w15_62),.acc(r15_62),.res(r15_63),.clk(clk),.wout(w15_63));
	PE pe15_64(.x(x64),.w(w15_63),.acc(r15_63),.res(r15_64),.clk(clk),.wout(w15_64));
	PE pe15_65(.x(x65),.w(w15_64),.acc(r15_64),.res(r15_65),.clk(clk),.wout(w15_65));
	PE pe15_66(.x(x66),.w(w15_65),.acc(r15_65),.res(r15_66),.clk(clk),.wout(w15_66));
	PE pe15_67(.x(x67),.w(w15_66),.acc(r15_66),.res(r15_67),.clk(clk),.wout(w15_67));
	PE pe15_68(.x(x68),.w(w15_67),.acc(r15_67),.res(r15_68),.clk(clk),.wout(w15_68));
	PE pe15_69(.x(x69),.w(w15_68),.acc(r15_68),.res(r15_69),.clk(clk),.wout(w15_69));
	PE pe15_70(.x(x70),.w(w15_69),.acc(r15_69),.res(r15_70),.clk(clk),.wout(w15_70));
	PE pe15_71(.x(x71),.w(w15_70),.acc(r15_70),.res(r15_71),.clk(clk),.wout(w15_71));
	PE pe15_72(.x(x72),.w(w15_71),.acc(r15_71),.res(r15_72),.clk(clk),.wout(w15_72));
	PE pe15_73(.x(x73),.w(w15_72),.acc(r15_72),.res(r15_73),.clk(clk),.wout(w15_73));
	PE pe15_74(.x(x74),.w(w15_73),.acc(r15_73),.res(r15_74),.clk(clk),.wout(w15_74));
	PE pe15_75(.x(x75),.w(w15_74),.acc(r15_74),.res(r15_75),.clk(clk),.wout(w15_75));
	PE pe15_76(.x(x76),.w(w15_75),.acc(r15_75),.res(r15_76),.clk(clk),.wout(w15_76));
	PE pe15_77(.x(x77),.w(w15_76),.acc(r15_76),.res(r15_77),.clk(clk),.wout(w15_77));
	PE pe15_78(.x(x78),.w(w15_77),.acc(r15_77),.res(r15_78),.clk(clk),.wout(w15_78));
	PE pe15_79(.x(x79),.w(w15_78),.acc(r15_78),.res(r15_79),.clk(clk),.wout(w15_79));
	PE pe15_80(.x(x80),.w(w15_79),.acc(r15_79),.res(r15_80),.clk(clk),.wout(w15_80));
	PE pe15_81(.x(x81),.w(w15_80),.acc(r15_80),.res(r15_81),.clk(clk),.wout(w15_81));
	PE pe15_82(.x(x82),.w(w15_81),.acc(r15_81),.res(r15_82),.clk(clk),.wout(w15_82));
	PE pe15_83(.x(x83),.w(w15_82),.acc(r15_82),.res(r15_83),.clk(clk),.wout(w15_83));
	PE pe15_84(.x(x84),.w(w15_83),.acc(r15_83),.res(r15_84),.clk(clk),.wout(w15_84));
	PE pe15_85(.x(x85),.w(w15_84),.acc(r15_84),.res(r15_85),.clk(clk),.wout(w15_85));
	PE pe15_86(.x(x86),.w(w15_85),.acc(r15_85),.res(r15_86),.clk(clk),.wout(w15_86));
	PE pe15_87(.x(x87),.w(w15_86),.acc(r15_86),.res(r15_87),.clk(clk),.wout(w15_87));
	PE pe15_88(.x(x88),.w(w15_87),.acc(r15_87),.res(r15_88),.clk(clk),.wout(w15_88));
	PE pe15_89(.x(x89),.w(w15_88),.acc(r15_88),.res(r15_89),.clk(clk),.wout(w15_89));
	PE pe15_90(.x(x90),.w(w15_89),.acc(r15_89),.res(r15_90),.clk(clk),.wout(w15_90));
	PE pe15_91(.x(x91),.w(w15_90),.acc(r15_90),.res(r15_91),.clk(clk),.wout(w15_91));
	PE pe15_92(.x(x92),.w(w15_91),.acc(r15_91),.res(r15_92),.clk(clk),.wout(w15_92));
	PE pe15_93(.x(x93),.w(w15_92),.acc(r15_92),.res(r15_93),.clk(clk),.wout(w15_93));
	PE pe15_94(.x(x94),.w(w15_93),.acc(r15_93),.res(r15_94),.clk(clk),.wout(w15_94));
	PE pe15_95(.x(x95),.w(w15_94),.acc(r15_94),.res(r15_95),.clk(clk),.wout(w15_95));
	PE pe15_96(.x(x96),.w(w15_95),.acc(r15_95),.res(r15_96),.clk(clk),.wout(w15_96));
	PE pe15_97(.x(x97),.w(w15_96),.acc(r15_96),.res(r15_97),.clk(clk),.wout(w15_97));
	PE pe15_98(.x(x98),.w(w15_97),.acc(r15_97),.res(r15_98),.clk(clk),.wout(w15_98));
	PE pe15_99(.x(x99),.w(w15_98),.acc(r15_98),.res(r15_99),.clk(clk),.wout(w15_99));
	PE pe15_100(.x(x100),.w(w15_99),.acc(r15_99),.res(r15_100),.clk(clk),.wout(w15_100));
	PE pe15_101(.x(x101),.w(w15_100),.acc(r15_100),.res(r15_101),.clk(clk),.wout(w15_101));
	PE pe15_102(.x(x102),.w(w15_101),.acc(r15_101),.res(r15_102),.clk(clk),.wout(w15_102));
	PE pe15_103(.x(x103),.w(w15_102),.acc(r15_102),.res(r15_103),.clk(clk),.wout(w15_103));
	PE pe15_104(.x(x104),.w(w15_103),.acc(r15_103),.res(r15_104),.clk(clk),.wout(w15_104));
	PE pe15_105(.x(x105),.w(w15_104),.acc(r15_104),.res(r15_105),.clk(clk),.wout(w15_105));
	PE pe15_106(.x(x106),.w(w15_105),.acc(r15_105),.res(r15_106),.clk(clk),.wout(w15_106));
	PE pe15_107(.x(x107),.w(w15_106),.acc(r15_106),.res(r15_107),.clk(clk),.wout(w15_107));
	PE pe15_108(.x(x108),.w(w15_107),.acc(r15_107),.res(r15_108),.clk(clk),.wout(w15_108));
	PE pe15_109(.x(x109),.w(w15_108),.acc(r15_108),.res(r15_109),.clk(clk),.wout(w15_109));
	PE pe15_110(.x(x110),.w(w15_109),.acc(r15_109),.res(r15_110),.clk(clk),.wout(w15_110));
	PE pe15_111(.x(x111),.w(w15_110),.acc(r15_110),.res(r15_111),.clk(clk),.wout(w15_111));
	PE pe15_112(.x(x112),.w(w15_111),.acc(r15_111),.res(r15_112),.clk(clk),.wout(w15_112));
	PE pe15_113(.x(x113),.w(w15_112),.acc(r15_112),.res(r15_113),.clk(clk),.wout(w15_113));
	PE pe15_114(.x(x114),.w(w15_113),.acc(r15_113),.res(r15_114),.clk(clk),.wout(w15_114));
	PE pe15_115(.x(x115),.w(w15_114),.acc(r15_114),.res(r15_115),.clk(clk),.wout(w15_115));
	PE pe15_116(.x(x116),.w(w15_115),.acc(r15_115),.res(r15_116),.clk(clk),.wout(w15_116));
	PE pe15_117(.x(x117),.w(w15_116),.acc(r15_116),.res(r15_117),.clk(clk),.wout(w15_117));
	PE pe15_118(.x(x118),.w(w15_117),.acc(r15_117),.res(r15_118),.clk(clk),.wout(w15_118));
	PE pe15_119(.x(x119),.w(w15_118),.acc(r15_118),.res(r15_119),.clk(clk),.wout(w15_119));
	PE pe15_120(.x(x120),.w(w15_119),.acc(r15_119),.res(r15_120),.clk(clk),.wout(w15_120));
	PE pe15_121(.x(x121),.w(w15_120),.acc(r15_120),.res(r15_121),.clk(clk),.wout(w15_121));
	PE pe15_122(.x(x122),.w(w15_121),.acc(r15_121),.res(r15_122),.clk(clk),.wout(w15_122));
	PE pe15_123(.x(x123),.w(w15_122),.acc(r15_122),.res(r15_123),.clk(clk),.wout(w15_123));
	PE pe15_124(.x(x124),.w(w15_123),.acc(r15_123),.res(r15_124),.clk(clk),.wout(w15_124));
	PE pe15_125(.x(x125),.w(w15_124),.acc(r15_124),.res(r15_125),.clk(clk),.wout(w15_125));
	PE pe15_126(.x(x126),.w(w15_125),.acc(r15_125),.res(r15_126),.clk(clk),.wout(w15_126));
	PE pe15_127(.x(x127),.w(w15_126),.acc(r15_126),.res(result15),.clk(clk),.wout(weight15));

	PE pe16_0(.x(x0),.w(w16),.acc(32'h0),.res(r16_0),.clk(clk),.wout(w16_0));
	PE pe16_1(.x(x1),.w(w16_0),.acc(r16_0),.res(r16_1),.clk(clk),.wout(w16_1));
	PE pe16_2(.x(x2),.w(w16_1),.acc(r16_1),.res(r16_2),.clk(clk),.wout(w16_2));
	PE pe16_3(.x(x3),.w(w16_2),.acc(r16_2),.res(r16_3),.clk(clk),.wout(w16_3));
	PE pe16_4(.x(x4),.w(w16_3),.acc(r16_3),.res(r16_4),.clk(clk),.wout(w16_4));
	PE pe16_5(.x(x5),.w(w16_4),.acc(r16_4),.res(r16_5),.clk(clk),.wout(w16_5));
	PE pe16_6(.x(x6),.w(w16_5),.acc(r16_5),.res(r16_6),.clk(clk),.wout(w16_6));
	PE pe16_7(.x(x7),.w(w16_6),.acc(r16_6),.res(r16_7),.clk(clk),.wout(w16_7));
	PE pe16_8(.x(x8),.w(w16_7),.acc(r16_7),.res(r16_8),.clk(clk),.wout(w16_8));
	PE pe16_9(.x(x9),.w(w16_8),.acc(r16_8),.res(r16_9),.clk(clk),.wout(w16_9));
	PE pe16_10(.x(x10),.w(w16_9),.acc(r16_9),.res(r16_10),.clk(clk),.wout(w16_10));
	PE pe16_11(.x(x11),.w(w16_10),.acc(r16_10),.res(r16_11),.clk(clk),.wout(w16_11));
	PE pe16_12(.x(x12),.w(w16_11),.acc(r16_11),.res(r16_12),.clk(clk),.wout(w16_12));
	PE pe16_13(.x(x13),.w(w16_12),.acc(r16_12),.res(r16_13),.clk(clk),.wout(w16_13));
	PE pe16_14(.x(x14),.w(w16_13),.acc(r16_13),.res(r16_14),.clk(clk),.wout(w16_14));
	PE pe16_15(.x(x15),.w(w16_14),.acc(r16_14),.res(r16_15),.clk(clk),.wout(w16_15));
	PE pe16_16(.x(x16),.w(w16_15),.acc(r16_15),.res(r16_16),.clk(clk),.wout(w16_16));
	PE pe16_17(.x(x17),.w(w16_16),.acc(r16_16),.res(r16_17),.clk(clk),.wout(w16_17));
	PE pe16_18(.x(x18),.w(w16_17),.acc(r16_17),.res(r16_18),.clk(clk),.wout(w16_18));
	PE pe16_19(.x(x19),.w(w16_18),.acc(r16_18),.res(r16_19),.clk(clk),.wout(w16_19));
	PE pe16_20(.x(x20),.w(w16_19),.acc(r16_19),.res(r16_20),.clk(clk),.wout(w16_20));
	PE pe16_21(.x(x21),.w(w16_20),.acc(r16_20),.res(r16_21),.clk(clk),.wout(w16_21));
	PE pe16_22(.x(x22),.w(w16_21),.acc(r16_21),.res(r16_22),.clk(clk),.wout(w16_22));
	PE pe16_23(.x(x23),.w(w16_22),.acc(r16_22),.res(r16_23),.clk(clk),.wout(w16_23));
	PE pe16_24(.x(x24),.w(w16_23),.acc(r16_23),.res(r16_24),.clk(clk),.wout(w16_24));
	PE pe16_25(.x(x25),.w(w16_24),.acc(r16_24),.res(r16_25),.clk(clk),.wout(w16_25));
	PE pe16_26(.x(x26),.w(w16_25),.acc(r16_25),.res(r16_26),.clk(clk),.wout(w16_26));
	PE pe16_27(.x(x27),.w(w16_26),.acc(r16_26),.res(r16_27),.clk(clk),.wout(w16_27));
	PE pe16_28(.x(x28),.w(w16_27),.acc(r16_27),.res(r16_28),.clk(clk),.wout(w16_28));
	PE pe16_29(.x(x29),.w(w16_28),.acc(r16_28),.res(r16_29),.clk(clk),.wout(w16_29));
	PE pe16_30(.x(x30),.w(w16_29),.acc(r16_29),.res(r16_30),.clk(clk),.wout(w16_30));
	PE pe16_31(.x(x31),.w(w16_30),.acc(r16_30),.res(r16_31),.clk(clk),.wout(w16_31));
	PE pe16_32(.x(x32),.w(w16_31),.acc(r16_31),.res(r16_32),.clk(clk),.wout(w16_32));
	PE pe16_33(.x(x33),.w(w16_32),.acc(r16_32),.res(r16_33),.clk(clk),.wout(w16_33));
	PE pe16_34(.x(x34),.w(w16_33),.acc(r16_33),.res(r16_34),.clk(clk),.wout(w16_34));
	PE pe16_35(.x(x35),.w(w16_34),.acc(r16_34),.res(r16_35),.clk(clk),.wout(w16_35));
	PE pe16_36(.x(x36),.w(w16_35),.acc(r16_35),.res(r16_36),.clk(clk),.wout(w16_36));
	PE pe16_37(.x(x37),.w(w16_36),.acc(r16_36),.res(r16_37),.clk(clk),.wout(w16_37));
	PE pe16_38(.x(x38),.w(w16_37),.acc(r16_37),.res(r16_38),.clk(clk),.wout(w16_38));
	PE pe16_39(.x(x39),.w(w16_38),.acc(r16_38),.res(r16_39),.clk(clk),.wout(w16_39));
	PE pe16_40(.x(x40),.w(w16_39),.acc(r16_39),.res(r16_40),.clk(clk),.wout(w16_40));
	PE pe16_41(.x(x41),.w(w16_40),.acc(r16_40),.res(r16_41),.clk(clk),.wout(w16_41));
	PE pe16_42(.x(x42),.w(w16_41),.acc(r16_41),.res(r16_42),.clk(clk),.wout(w16_42));
	PE pe16_43(.x(x43),.w(w16_42),.acc(r16_42),.res(r16_43),.clk(clk),.wout(w16_43));
	PE pe16_44(.x(x44),.w(w16_43),.acc(r16_43),.res(r16_44),.clk(clk),.wout(w16_44));
	PE pe16_45(.x(x45),.w(w16_44),.acc(r16_44),.res(r16_45),.clk(clk),.wout(w16_45));
	PE pe16_46(.x(x46),.w(w16_45),.acc(r16_45),.res(r16_46),.clk(clk),.wout(w16_46));
	PE pe16_47(.x(x47),.w(w16_46),.acc(r16_46),.res(r16_47),.clk(clk),.wout(w16_47));
	PE pe16_48(.x(x48),.w(w16_47),.acc(r16_47),.res(r16_48),.clk(clk),.wout(w16_48));
	PE pe16_49(.x(x49),.w(w16_48),.acc(r16_48),.res(r16_49),.clk(clk),.wout(w16_49));
	PE pe16_50(.x(x50),.w(w16_49),.acc(r16_49),.res(r16_50),.clk(clk),.wout(w16_50));
	PE pe16_51(.x(x51),.w(w16_50),.acc(r16_50),.res(r16_51),.clk(clk),.wout(w16_51));
	PE pe16_52(.x(x52),.w(w16_51),.acc(r16_51),.res(r16_52),.clk(clk),.wout(w16_52));
	PE pe16_53(.x(x53),.w(w16_52),.acc(r16_52),.res(r16_53),.clk(clk),.wout(w16_53));
	PE pe16_54(.x(x54),.w(w16_53),.acc(r16_53),.res(r16_54),.clk(clk),.wout(w16_54));
	PE pe16_55(.x(x55),.w(w16_54),.acc(r16_54),.res(r16_55),.clk(clk),.wout(w16_55));
	PE pe16_56(.x(x56),.w(w16_55),.acc(r16_55),.res(r16_56),.clk(clk),.wout(w16_56));
	PE pe16_57(.x(x57),.w(w16_56),.acc(r16_56),.res(r16_57),.clk(clk),.wout(w16_57));
	PE pe16_58(.x(x58),.w(w16_57),.acc(r16_57),.res(r16_58),.clk(clk),.wout(w16_58));
	PE pe16_59(.x(x59),.w(w16_58),.acc(r16_58),.res(r16_59),.clk(clk),.wout(w16_59));
	PE pe16_60(.x(x60),.w(w16_59),.acc(r16_59),.res(r16_60),.clk(clk),.wout(w16_60));
	PE pe16_61(.x(x61),.w(w16_60),.acc(r16_60),.res(r16_61),.clk(clk),.wout(w16_61));
	PE pe16_62(.x(x62),.w(w16_61),.acc(r16_61),.res(r16_62),.clk(clk),.wout(w16_62));
	PE pe16_63(.x(x63),.w(w16_62),.acc(r16_62),.res(r16_63),.clk(clk),.wout(w16_63));
	PE pe16_64(.x(x64),.w(w16_63),.acc(r16_63),.res(r16_64),.clk(clk),.wout(w16_64));
	PE pe16_65(.x(x65),.w(w16_64),.acc(r16_64),.res(r16_65),.clk(clk),.wout(w16_65));
	PE pe16_66(.x(x66),.w(w16_65),.acc(r16_65),.res(r16_66),.clk(clk),.wout(w16_66));
	PE pe16_67(.x(x67),.w(w16_66),.acc(r16_66),.res(r16_67),.clk(clk),.wout(w16_67));
	PE pe16_68(.x(x68),.w(w16_67),.acc(r16_67),.res(r16_68),.clk(clk),.wout(w16_68));
	PE pe16_69(.x(x69),.w(w16_68),.acc(r16_68),.res(r16_69),.clk(clk),.wout(w16_69));
	PE pe16_70(.x(x70),.w(w16_69),.acc(r16_69),.res(r16_70),.clk(clk),.wout(w16_70));
	PE pe16_71(.x(x71),.w(w16_70),.acc(r16_70),.res(r16_71),.clk(clk),.wout(w16_71));
	PE pe16_72(.x(x72),.w(w16_71),.acc(r16_71),.res(r16_72),.clk(clk),.wout(w16_72));
	PE pe16_73(.x(x73),.w(w16_72),.acc(r16_72),.res(r16_73),.clk(clk),.wout(w16_73));
	PE pe16_74(.x(x74),.w(w16_73),.acc(r16_73),.res(r16_74),.clk(clk),.wout(w16_74));
	PE pe16_75(.x(x75),.w(w16_74),.acc(r16_74),.res(r16_75),.clk(clk),.wout(w16_75));
	PE pe16_76(.x(x76),.w(w16_75),.acc(r16_75),.res(r16_76),.clk(clk),.wout(w16_76));
	PE pe16_77(.x(x77),.w(w16_76),.acc(r16_76),.res(r16_77),.clk(clk),.wout(w16_77));
	PE pe16_78(.x(x78),.w(w16_77),.acc(r16_77),.res(r16_78),.clk(clk),.wout(w16_78));
	PE pe16_79(.x(x79),.w(w16_78),.acc(r16_78),.res(r16_79),.clk(clk),.wout(w16_79));
	PE pe16_80(.x(x80),.w(w16_79),.acc(r16_79),.res(r16_80),.clk(clk),.wout(w16_80));
	PE pe16_81(.x(x81),.w(w16_80),.acc(r16_80),.res(r16_81),.clk(clk),.wout(w16_81));
	PE pe16_82(.x(x82),.w(w16_81),.acc(r16_81),.res(r16_82),.clk(clk),.wout(w16_82));
	PE pe16_83(.x(x83),.w(w16_82),.acc(r16_82),.res(r16_83),.clk(clk),.wout(w16_83));
	PE pe16_84(.x(x84),.w(w16_83),.acc(r16_83),.res(r16_84),.clk(clk),.wout(w16_84));
	PE pe16_85(.x(x85),.w(w16_84),.acc(r16_84),.res(r16_85),.clk(clk),.wout(w16_85));
	PE pe16_86(.x(x86),.w(w16_85),.acc(r16_85),.res(r16_86),.clk(clk),.wout(w16_86));
	PE pe16_87(.x(x87),.w(w16_86),.acc(r16_86),.res(r16_87),.clk(clk),.wout(w16_87));
	PE pe16_88(.x(x88),.w(w16_87),.acc(r16_87),.res(r16_88),.clk(clk),.wout(w16_88));
	PE pe16_89(.x(x89),.w(w16_88),.acc(r16_88),.res(r16_89),.clk(clk),.wout(w16_89));
	PE pe16_90(.x(x90),.w(w16_89),.acc(r16_89),.res(r16_90),.clk(clk),.wout(w16_90));
	PE pe16_91(.x(x91),.w(w16_90),.acc(r16_90),.res(r16_91),.clk(clk),.wout(w16_91));
	PE pe16_92(.x(x92),.w(w16_91),.acc(r16_91),.res(r16_92),.clk(clk),.wout(w16_92));
	PE pe16_93(.x(x93),.w(w16_92),.acc(r16_92),.res(r16_93),.clk(clk),.wout(w16_93));
	PE pe16_94(.x(x94),.w(w16_93),.acc(r16_93),.res(r16_94),.clk(clk),.wout(w16_94));
	PE pe16_95(.x(x95),.w(w16_94),.acc(r16_94),.res(r16_95),.clk(clk),.wout(w16_95));
	PE pe16_96(.x(x96),.w(w16_95),.acc(r16_95),.res(r16_96),.clk(clk),.wout(w16_96));
	PE pe16_97(.x(x97),.w(w16_96),.acc(r16_96),.res(r16_97),.clk(clk),.wout(w16_97));
	PE pe16_98(.x(x98),.w(w16_97),.acc(r16_97),.res(r16_98),.clk(clk),.wout(w16_98));
	PE pe16_99(.x(x99),.w(w16_98),.acc(r16_98),.res(r16_99),.clk(clk),.wout(w16_99));
	PE pe16_100(.x(x100),.w(w16_99),.acc(r16_99),.res(r16_100),.clk(clk),.wout(w16_100));
	PE pe16_101(.x(x101),.w(w16_100),.acc(r16_100),.res(r16_101),.clk(clk),.wout(w16_101));
	PE pe16_102(.x(x102),.w(w16_101),.acc(r16_101),.res(r16_102),.clk(clk),.wout(w16_102));
	PE pe16_103(.x(x103),.w(w16_102),.acc(r16_102),.res(r16_103),.clk(clk),.wout(w16_103));
	PE pe16_104(.x(x104),.w(w16_103),.acc(r16_103),.res(r16_104),.clk(clk),.wout(w16_104));
	PE pe16_105(.x(x105),.w(w16_104),.acc(r16_104),.res(r16_105),.clk(clk),.wout(w16_105));
	PE pe16_106(.x(x106),.w(w16_105),.acc(r16_105),.res(r16_106),.clk(clk),.wout(w16_106));
	PE pe16_107(.x(x107),.w(w16_106),.acc(r16_106),.res(r16_107),.clk(clk),.wout(w16_107));
	PE pe16_108(.x(x108),.w(w16_107),.acc(r16_107),.res(r16_108),.clk(clk),.wout(w16_108));
	PE pe16_109(.x(x109),.w(w16_108),.acc(r16_108),.res(r16_109),.clk(clk),.wout(w16_109));
	PE pe16_110(.x(x110),.w(w16_109),.acc(r16_109),.res(r16_110),.clk(clk),.wout(w16_110));
	PE pe16_111(.x(x111),.w(w16_110),.acc(r16_110),.res(r16_111),.clk(clk),.wout(w16_111));
	PE pe16_112(.x(x112),.w(w16_111),.acc(r16_111),.res(r16_112),.clk(clk),.wout(w16_112));
	PE pe16_113(.x(x113),.w(w16_112),.acc(r16_112),.res(r16_113),.clk(clk),.wout(w16_113));
	PE pe16_114(.x(x114),.w(w16_113),.acc(r16_113),.res(r16_114),.clk(clk),.wout(w16_114));
	PE pe16_115(.x(x115),.w(w16_114),.acc(r16_114),.res(r16_115),.clk(clk),.wout(w16_115));
	PE pe16_116(.x(x116),.w(w16_115),.acc(r16_115),.res(r16_116),.clk(clk),.wout(w16_116));
	PE pe16_117(.x(x117),.w(w16_116),.acc(r16_116),.res(r16_117),.clk(clk),.wout(w16_117));
	PE pe16_118(.x(x118),.w(w16_117),.acc(r16_117),.res(r16_118),.clk(clk),.wout(w16_118));
	PE pe16_119(.x(x119),.w(w16_118),.acc(r16_118),.res(r16_119),.clk(clk),.wout(w16_119));
	PE pe16_120(.x(x120),.w(w16_119),.acc(r16_119),.res(r16_120),.clk(clk),.wout(w16_120));
	PE pe16_121(.x(x121),.w(w16_120),.acc(r16_120),.res(r16_121),.clk(clk),.wout(w16_121));
	PE pe16_122(.x(x122),.w(w16_121),.acc(r16_121),.res(r16_122),.clk(clk),.wout(w16_122));
	PE pe16_123(.x(x123),.w(w16_122),.acc(r16_122),.res(r16_123),.clk(clk),.wout(w16_123));
	PE pe16_124(.x(x124),.w(w16_123),.acc(r16_123),.res(r16_124),.clk(clk),.wout(w16_124));
	PE pe16_125(.x(x125),.w(w16_124),.acc(r16_124),.res(r16_125),.clk(clk),.wout(w16_125));
	PE pe16_126(.x(x126),.w(w16_125),.acc(r16_125),.res(r16_126),.clk(clk),.wout(w16_126));
	PE pe16_127(.x(x127),.w(w16_126),.acc(r16_126),.res(result16),.clk(clk),.wout(weight16));

	PE pe17_0(.x(x0),.w(w17),.acc(32'h0),.res(r17_0),.clk(clk),.wout(w17_0));
	PE pe17_1(.x(x1),.w(w17_0),.acc(r17_0),.res(r17_1),.clk(clk),.wout(w17_1));
	PE pe17_2(.x(x2),.w(w17_1),.acc(r17_1),.res(r17_2),.clk(clk),.wout(w17_2));
	PE pe17_3(.x(x3),.w(w17_2),.acc(r17_2),.res(r17_3),.clk(clk),.wout(w17_3));
	PE pe17_4(.x(x4),.w(w17_3),.acc(r17_3),.res(r17_4),.clk(clk),.wout(w17_4));
	PE pe17_5(.x(x5),.w(w17_4),.acc(r17_4),.res(r17_5),.clk(clk),.wout(w17_5));
	PE pe17_6(.x(x6),.w(w17_5),.acc(r17_5),.res(r17_6),.clk(clk),.wout(w17_6));
	PE pe17_7(.x(x7),.w(w17_6),.acc(r17_6),.res(r17_7),.clk(clk),.wout(w17_7));
	PE pe17_8(.x(x8),.w(w17_7),.acc(r17_7),.res(r17_8),.clk(clk),.wout(w17_8));
	PE pe17_9(.x(x9),.w(w17_8),.acc(r17_8),.res(r17_9),.clk(clk),.wout(w17_9));
	PE pe17_10(.x(x10),.w(w17_9),.acc(r17_9),.res(r17_10),.clk(clk),.wout(w17_10));
	PE pe17_11(.x(x11),.w(w17_10),.acc(r17_10),.res(r17_11),.clk(clk),.wout(w17_11));
	PE pe17_12(.x(x12),.w(w17_11),.acc(r17_11),.res(r17_12),.clk(clk),.wout(w17_12));
	PE pe17_13(.x(x13),.w(w17_12),.acc(r17_12),.res(r17_13),.clk(clk),.wout(w17_13));
	PE pe17_14(.x(x14),.w(w17_13),.acc(r17_13),.res(r17_14),.clk(clk),.wout(w17_14));
	PE pe17_15(.x(x15),.w(w17_14),.acc(r17_14),.res(r17_15),.clk(clk),.wout(w17_15));
	PE pe17_16(.x(x16),.w(w17_15),.acc(r17_15),.res(r17_16),.clk(clk),.wout(w17_16));
	PE pe17_17(.x(x17),.w(w17_16),.acc(r17_16),.res(r17_17),.clk(clk),.wout(w17_17));
	PE pe17_18(.x(x18),.w(w17_17),.acc(r17_17),.res(r17_18),.clk(clk),.wout(w17_18));
	PE pe17_19(.x(x19),.w(w17_18),.acc(r17_18),.res(r17_19),.clk(clk),.wout(w17_19));
	PE pe17_20(.x(x20),.w(w17_19),.acc(r17_19),.res(r17_20),.clk(clk),.wout(w17_20));
	PE pe17_21(.x(x21),.w(w17_20),.acc(r17_20),.res(r17_21),.clk(clk),.wout(w17_21));
	PE pe17_22(.x(x22),.w(w17_21),.acc(r17_21),.res(r17_22),.clk(clk),.wout(w17_22));
	PE pe17_23(.x(x23),.w(w17_22),.acc(r17_22),.res(r17_23),.clk(clk),.wout(w17_23));
	PE pe17_24(.x(x24),.w(w17_23),.acc(r17_23),.res(r17_24),.clk(clk),.wout(w17_24));
	PE pe17_25(.x(x25),.w(w17_24),.acc(r17_24),.res(r17_25),.clk(clk),.wout(w17_25));
	PE pe17_26(.x(x26),.w(w17_25),.acc(r17_25),.res(r17_26),.clk(clk),.wout(w17_26));
	PE pe17_27(.x(x27),.w(w17_26),.acc(r17_26),.res(r17_27),.clk(clk),.wout(w17_27));
	PE pe17_28(.x(x28),.w(w17_27),.acc(r17_27),.res(r17_28),.clk(clk),.wout(w17_28));
	PE pe17_29(.x(x29),.w(w17_28),.acc(r17_28),.res(r17_29),.clk(clk),.wout(w17_29));
	PE pe17_30(.x(x30),.w(w17_29),.acc(r17_29),.res(r17_30),.clk(clk),.wout(w17_30));
	PE pe17_31(.x(x31),.w(w17_30),.acc(r17_30),.res(r17_31),.clk(clk),.wout(w17_31));
	PE pe17_32(.x(x32),.w(w17_31),.acc(r17_31),.res(r17_32),.clk(clk),.wout(w17_32));
	PE pe17_33(.x(x33),.w(w17_32),.acc(r17_32),.res(r17_33),.clk(clk),.wout(w17_33));
	PE pe17_34(.x(x34),.w(w17_33),.acc(r17_33),.res(r17_34),.clk(clk),.wout(w17_34));
	PE pe17_35(.x(x35),.w(w17_34),.acc(r17_34),.res(r17_35),.clk(clk),.wout(w17_35));
	PE pe17_36(.x(x36),.w(w17_35),.acc(r17_35),.res(r17_36),.clk(clk),.wout(w17_36));
	PE pe17_37(.x(x37),.w(w17_36),.acc(r17_36),.res(r17_37),.clk(clk),.wout(w17_37));
	PE pe17_38(.x(x38),.w(w17_37),.acc(r17_37),.res(r17_38),.clk(clk),.wout(w17_38));
	PE pe17_39(.x(x39),.w(w17_38),.acc(r17_38),.res(r17_39),.clk(clk),.wout(w17_39));
	PE pe17_40(.x(x40),.w(w17_39),.acc(r17_39),.res(r17_40),.clk(clk),.wout(w17_40));
	PE pe17_41(.x(x41),.w(w17_40),.acc(r17_40),.res(r17_41),.clk(clk),.wout(w17_41));
	PE pe17_42(.x(x42),.w(w17_41),.acc(r17_41),.res(r17_42),.clk(clk),.wout(w17_42));
	PE pe17_43(.x(x43),.w(w17_42),.acc(r17_42),.res(r17_43),.clk(clk),.wout(w17_43));
	PE pe17_44(.x(x44),.w(w17_43),.acc(r17_43),.res(r17_44),.clk(clk),.wout(w17_44));
	PE pe17_45(.x(x45),.w(w17_44),.acc(r17_44),.res(r17_45),.clk(clk),.wout(w17_45));
	PE pe17_46(.x(x46),.w(w17_45),.acc(r17_45),.res(r17_46),.clk(clk),.wout(w17_46));
	PE pe17_47(.x(x47),.w(w17_46),.acc(r17_46),.res(r17_47),.clk(clk),.wout(w17_47));
	PE pe17_48(.x(x48),.w(w17_47),.acc(r17_47),.res(r17_48),.clk(clk),.wout(w17_48));
	PE pe17_49(.x(x49),.w(w17_48),.acc(r17_48),.res(r17_49),.clk(clk),.wout(w17_49));
	PE pe17_50(.x(x50),.w(w17_49),.acc(r17_49),.res(r17_50),.clk(clk),.wout(w17_50));
	PE pe17_51(.x(x51),.w(w17_50),.acc(r17_50),.res(r17_51),.clk(clk),.wout(w17_51));
	PE pe17_52(.x(x52),.w(w17_51),.acc(r17_51),.res(r17_52),.clk(clk),.wout(w17_52));
	PE pe17_53(.x(x53),.w(w17_52),.acc(r17_52),.res(r17_53),.clk(clk),.wout(w17_53));
	PE pe17_54(.x(x54),.w(w17_53),.acc(r17_53),.res(r17_54),.clk(clk),.wout(w17_54));
	PE pe17_55(.x(x55),.w(w17_54),.acc(r17_54),.res(r17_55),.clk(clk),.wout(w17_55));
	PE pe17_56(.x(x56),.w(w17_55),.acc(r17_55),.res(r17_56),.clk(clk),.wout(w17_56));
	PE pe17_57(.x(x57),.w(w17_56),.acc(r17_56),.res(r17_57),.clk(clk),.wout(w17_57));
	PE pe17_58(.x(x58),.w(w17_57),.acc(r17_57),.res(r17_58),.clk(clk),.wout(w17_58));
	PE pe17_59(.x(x59),.w(w17_58),.acc(r17_58),.res(r17_59),.clk(clk),.wout(w17_59));
	PE pe17_60(.x(x60),.w(w17_59),.acc(r17_59),.res(r17_60),.clk(clk),.wout(w17_60));
	PE pe17_61(.x(x61),.w(w17_60),.acc(r17_60),.res(r17_61),.clk(clk),.wout(w17_61));
	PE pe17_62(.x(x62),.w(w17_61),.acc(r17_61),.res(r17_62),.clk(clk),.wout(w17_62));
	PE pe17_63(.x(x63),.w(w17_62),.acc(r17_62),.res(r17_63),.clk(clk),.wout(w17_63));
	PE pe17_64(.x(x64),.w(w17_63),.acc(r17_63),.res(r17_64),.clk(clk),.wout(w17_64));
	PE pe17_65(.x(x65),.w(w17_64),.acc(r17_64),.res(r17_65),.clk(clk),.wout(w17_65));
	PE pe17_66(.x(x66),.w(w17_65),.acc(r17_65),.res(r17_66),.clk(clk),.wout(w17_66));
	PE pe17_67(.x(x67),.w(w17_66),.acc(r17_66),.res(r17_67),.clk(clk),.wout(w17_67));
	PE pe17_68(.x(x68),.w(w17_67),.acc(r17_67),.res(r17_68),.clk(clk),.wout(w17_68));
	PE pe17_69(.x(x69),.w(w17_68),.acc(r17_68),.res(r17_69),.clk(clk),.wout(w17_69));
	PE pe17_70(.x(x70),.w(w17_69),.acc(r17_69),.res(r17_70),.clk(clk),.wout(w17_70));
	PE pe17_71(.x(x71),.w(w17_70),.acc(r17_70),.res(r17_71),.clk(clk),.wout(w17_71));
	PE pe17_72(.x(x72),.w(w17_71),.acc(r17_71),.res(r17_72),.clk(clk),.wout(w17_72));
	PE pe17_73(.x(x73),.w(w17_72),.acc(r17_72),.res(r17_73),.clk(clk),.wout(w17_73));
	PE pe17_74(.x(x74),.w(w17_73),.acc(r17_73),.res(r17_74),.clk(clk),.wout(w17_74));
	PE pe17_75(.x(x75),.w(w17_74),.acc(r17_74),.res(r17_75),.clk(clk),.wout(w17_75));
	PE pe17_76(.x(x76),.w(w17_75),.acc(r17_75),.res(r17_76),.clk(clk),.wout(w17_76));
	PE pe17_77(.x(x77),.w(w17_76),.acc(r17_76),.res(r17_77),.clk(clk),.wout(w17_77));
	PE pe17_78(.x(x78),.w(w17_77),.acc(r17_77),.res(r17_78),.clk(clk),.wout(w17_78));
	PE pe17_79(.x(x79),.w(w17_78),.acc(r17_78),.res(r17_79),.clk(clk),.wout(w17_79));
	PE pe17_80(.x(x80),.w(w17_79),.acc(r17_79),.res(r17_80),.clk(clk),.wout(w17_80));
	PE pe17_81(.x(x81),.w(w17_80),.acc(r17_80),.res(r17_81),.clk(clk),.wout(w17_81));
	PE pe17_82(.x(x82),.w(w17_81),.acc(r17_81),.res(r17_82),.clk(clk),.wout(w17_82));
	PE pe17_83(.x(x83),.w(w17_82),.acc(r17_82),.res(r17_83),.clk(clk),.wout(w17_83));
	PE pe17_84(.x(x84),.w(w17_83),.acc(r17_83),.res(r17_84),.clk(clk),.wout(w17_84));
	PE pe17_85(.x(x85),.w(w17_84),.acc(r17_84),.res(r17_85),.clk(clk),.wout(w17_85));
	PE pe17_86(.x(x86),.w(w17_85),.acc(r17_85),.res(r17_86),.clk(clk),.wout(w17_86));
	PE pe17_87(.x(x87),.w(w17_86),.acc(r17_86),.res(r17_87),.clk(clk),.wout(w17_87));
	PE pe17_88(.x(x88),.w(w17_87),.acc(r17_87),.res(r17_88),.clk(clk),.wout(w17_88));
	PE pe17_89(.x(x89),.w(w17_88),.acc(r17_88),.res(r17_89),.clk(clk),.wout(w17_89));
	PE pe17_90(.x(x90),.w(w17_89),.acc(r17_89),.res(r17_90),.clk(clk),.wout(w17_90));
	PE pe17_91(.x(x91),.w(w17_90),.acc(r17_90),.res(r17_91),.clk(clk),.wout(w17_91));
	PE pe17_92(.x(x92),.w(w17_91),.acc(r17_91),.res(r17_92),.clk(clk),.wout(w17_92));
	PE pe17_93(.x(x93),.w(w17_92),.acc(r17_92),.res(r17_93),.clk(clk),.wout(w17_93));
	PE pe17_94(.x(x94),.w(w17_93),.acc(r17_93),.res(r17_94),.clk(clk),.wout(w17_94));
	PE pe17_95(.x(x95),.w(w17_94),.acc(r17_94),.res(r17_95),.clk(clk),.wout(w17_95));
	PE pe17_96(.x(x96),.w(w17_95),.acc(r17_95),.res(r17_96),.clk(clk),.wout(w17_96));
	PE pe17_97(.x(x97),.w(w17_96),.acc(r17_96),.res(r17_97),.clk(clk),.wout(w17_97));
	PE pe17_98(.x(x98),.w(w17_97),.acc(r17_97),.res(r17_98),.clk(clk),.wout(w17_98));
	PE pe17_99(.x(x99),.w(w17_98),.acc(r17_98),.res(r17_99),.clk(clk),.wout(w17_99));
	PE pe17_100(.x(x100),.w(w17_99),.acc(r17_99),.res(r17_100),.clk(clk),.wout(w17_100));
	PE pe17_101(.x(x101),.w(w17_100),.acc(r17_100),.res(r17_101),.clk(clk),.wout(w17_101));
	PE pe17_102(.x(x102),.w(w17_101),.acc(r17_101),.res(r17_102),.clk(clk),.wout(w17_102));
	PE pe17_103(.x(x103),.w(w17_102),.acc(r17_102),.res(r17_103),.clk(clk),.wout(w17_103));
	PE pe17_104(.x(x104),.w(w17_103),.acc(r17_103),.res(r17_104),.clk(clk),.wout(w17_104));
	PE pe17_105(.x(x105),.w(w17_104),.acc(r17_104),.res(r17_105),.clk(clk),.wout(w17_105));
	PE pe17_106(.x(x106),.w(w17_105),.acc(r17_105),.res(r17_106),.clk(clk),.wout(w17_106));
	PE pe17_107(.x(x107),.w(w17_106),.acc(r17_106),.res(r17_107),.clk(clk),.wout(w17_107));
	PE pe17_108(.x(x108),.w(w17_107),.acc(r17_107),.res(r17_108),.clk(clk),.wout(w17_108));
	PE pe17_109(.x(x109),.w(w17_108),.acc(r17_108),.res(r17_109),.clk(clk),.wout(w17_109));
	PE pe17_110(.x(x110),.w(w17_109),.acc(r17_109),.res(r17_110),.clk(clk),.wout(w17_110));
	PE pe17_111(.x(x111),.w(w17_110),.acc(r17_110),.res(r17_111),.clk(clk),.wout(w17_111));
	PE pe17_112(.x(x112),.w(w17_111),.acc(r17_111),.res(r17_112),.clk(clk),.wout(w17_112));
	PE pe17_113(.x(x113),.w(w17_112),.acc(r17_112),.res(r17_113),.clk(clk),.wout(w17_113));
	PE pe17_114(.x(x114),.w(w17_113),.acc(r17_113),.res(r17_114),.clk(clk),.wout(w17_114));
	PE pe17_115(.x(x115),.w(w17_114),.acc(r17_114),.res(r17_115),.clk(clk),.wout(w17_115));
	PE pe17_116(.x(x116),.w(w17_115),.acc(r17_115),.res(r17_116),.clk(clk),.wout(w17_116));
	PE pe17_117(.x(x117),.w(w17_116),.acc(r17_116),.res(r17_117),.clk(clk),.wout(w17_117));
	PE pe17_118(.x(x118),.w(w17_117),.acc(r17_117),.res(r17_118),.clk(clk),.wout(w17_118));
	PE pe17_119(.x(x119),.w(w17_118),.acc(r17_118),.res(r17_119),.clk(clk),.wout(w17_119));
	PE pe17_120(.x(x120),.w(w17_119),.acc(r17_119),.res(r17_120),.clk(clk),.wout(w17_120));
	PE pe17_121(.x(x121),.w(w17_120),.acc(r17_120),.res(r17_121),.clk(clk),.wout(w17_121));
	PE pe17_122(.x(x122),.w(w17_121),.acc(r17_121),.res(r17_122),.clk(clk),.wout(w17_122));
	PE pe17_123(.x(x123),.w(w17_122),.acc(r17_122),.res(r17_123),.clk(clk),.wout(w17_123));
	PE pe17_124(.x(x124),.w(w17_123),.acc(r17_123),.res(r17_124),.clk(clk),.wout(w17_124));
	PE pe17_125(.x(x125),.w(w17_124),.acc(r17_124),.res(r17_125),.clk(clk),.wout(w17_125));
	PE pe17_126(.x(x126),.w(w17_125),.acc(r17_125),.res(r17_126),.clk(clk),.wout(w17_126));
	PE pe17_127(.x(x127),.w(w17_126),.acc(r17_126),.res(result17),.clk(clk),.wout(weight17));

	PE pe18_0(.x(x0),.w(w18),.acc(32'h0),.res(r18_0),.clk(clk),.wout(w18_0));
	PE pe18_1(.x(x1),.w(w18_0),.acc(r18_0),.res(r18_1),.clk(clk),.wout(w18_1));
	PE pe18_2(.x(x2),.w(w18_1),.acc(r18_1),.res(r18_2),.clk(clk),.wout(w18_2));
	PE pe18_3(.x(x3),.w(w18_2),.acc(r18_2),.res(r18_3),.clk(clk),.wout(w18_3));
	PE pe18_4(.x(x4),.w(w18_3),.acc(r18_3),.res(r18_4),.clk(clk),.wout(w18_4));
	PE pe18_5(.x(x5),.w(w18_4),.acc(r18_4),.res(r18_5),.clk(clk),.wout(w18_5));
	PE pe18_6(.x(x6),.w(w18_5),.acc(r18_5),.res(r18_6),.clk(clk),.wout(w18_6));
	PE pe18_7(.x(x7),.w(w18_6),.acc(r18_6),.res(r18_7),.clk(clk),.wout(w18_7));
	PE pe18_8(.x(x8),.w(w18_7),.acc(r18_7),.res(r18_8),.clk(clk),.wout(w18_8));
	PE pe18_9(.x(x9),.w(w18_8),.acc(r18_8),.res(r18_9),.clk(clk),.wout(w18_9));
	PE pe18_10(.x(x10),.w(w18_9),.acc(r18_9),.res(r18_10),.clk(clk),.wout(w18_10));
	PE pe18_11(.x(x11),.w(w18_10),.acc(r18_10),.res(r18_11),.clk(clk),.wout(w18_11));
	PE pe18_12(.x(x12),.w(w18_11),.acc(r18_11),.res(r18_12),.clk(clk),.wout(w18_12));
	PE pe18_13(.x(x13),.w(w18_12),.acc(r18_12),.res(r18_13),.clk(clk),.wout(w18_13));
	PE pe18_14(.x(x14),.w(w18_13),.acc(r18_13),.res(r18_14),.clk(clk),.wout(w18_14));
	PE pe18_15(.x(x15),.w(w18_14),.acc(r18_14),.res(r18_15),.clk(clk),.wout(w18_15));
	PE pe18_16(.x(x16),.w(w18_15),.acc(r18_15),.res(r18_16),.clk(clk),.wout(w18_16));
	PE pe18_17(.x(x17),.w(w18_16),.acc(r18_16),.res(r18_17),.clk(clk),.wout(w18_17));
	PE pe18_18(.x(x18),.w(w18_17),.acc(r18_17),.res(r18_18),.clk(clk),.wout(w18_18));
	PE pe18_19(.x(x19),.w(w18_18),.acc(r18_18),.res(r18_19),.clk(clk),.wout(w18_19));
	PE pe18_20(.x(x20),.w(w18_19),.acc(r18_19),.res(r18_20),.clk(clk),.wout(w18_20));
	PE pe18_21(.x(x21),.w(w18_20),.acc(r18_20),.res(r18_21),.clk(clk),.wout(w18_21));
	PE pe18_22(.x(x22),.w(w18_21),.acc(r18_21),.res(r18_22),.clk(clk),.wout(w18_22));
	PE pe18_23(.x(x23),.w(w18_22),.acc(r18_22),.res(r18_23),.clk(clk),.wout(w18_23));
	PE pe18_24(.x(x24),.w(w18_23),.acc(r18_23),.res(r18_24),.clk(clk),.wout(w18_24));
	PE pe18_25(.x(x25),.w(w18_24),.acc(r18_24),.res(r18_25),.clk(clk),.wout(w18_25));
	PE pe18_26(.x(x26),.w(w18_25),.acc(r18_25),.res(r18_26),.clk(clk),.wout(w18_26));
	PE pe18_27(.x(x27),.w(w18_26),.acc(r18_26),.res(r18_27),.clk(clk),.wout(w18_27));
	PE pe18_28(.x(x28),.w(w18_27),.acc(r18_27),.res(r18_28),.clk(clk),.wout(w18_28));
	PE pe18_29(.x(x29),.w(w18_28),.acc(r18_28),.res(r18_29),.clk(clk),.wout(w18_29));
	PE pe18_30(.x(x30),.w(w18_29),.acc(r18_29),.res(r18_30),.clk(clk),.wout(w18_30));
	PE pe18_31(.x(x31),.w(w18_30),.acc(r18_30),.res(r18_31),.clk(clk),.wout(w18_31));
	PE pe18_32(.x(x32),.w(w18_31),.acc(r18_31),.res(r18_32),.clk(clk),.wout(w18_32));
	PE pe18_33(.x(x33),.w(w18_32),.acc(r18_32),.res(r18_33),.clk(clk),.wout(w18_33));
	PE pe18_34(.x(x34),.w(w18_33),.acc(r18_33),.res(r18_34),.clk(clk),.wout(w18_34));
	PE pe18_35(.x(x35),.w(w18_34),.acc(r18_34),.res(r18_35),.clk(clk),.wout(w18_35));
	PE pe18_36(.x(x36),.w(w18_35),.acc(r18_35),.res(r18_36),.clk(clk),.wout(w18_36));
	PE pe18_37(.x(x37),.w(w18_36),.acc(r18_36),.res(r18_37),.clk(clk),.wout(w18_37));
	PE pe18_38(.x(x38),.w(w18_37),.acc(r18_37),.res(r18_38),.clk(clk),.wout(w18_38));
	PE pe18_39(.x(x39),.w(w18_38),.acc(r18_38),.res(r18_39),.clk(clk),.wout(w18_39));
	PE pe18_40(.x(x40),.w(w18_39),.acc(r18_39),.res(r18_40),.clk(clk),.wout(w18_40));
	PE pe18_41(.x(x41),.w(w18_40),.acc(r18_40),.res(r18_41),.clk(clk),.wout(w18_41));
	PE pe18_42(.x(x42),.w(w18_41),.acc(r18_41),.res(r18_42),.clk(clk),.wout(w18_42));
	PE pe18_43(.x(x43),.w(w18_42),.acc(r18_42),.res(r18_43),.clk(clk),.wout(w18_43));
	PE pe18_44(.x(x44),.w(w18_43),.acc(r18_43),.res(r18_44),.clk(clk),.wout(w18_44));
	PE pe18_45(.x(x45),.w(w18_44),.acc(r18_44),.res(r18_45),.clk(clk),.wout(w18_45));
	PE pe18_46(.x(x46),.w(w18_45),.acc(r18_45),.res(r18_46),.clk(clk),.wout(w18_46));
	PE pe18_47(.x(x47),.w(w18_46),.acc(r18_46),.res(r18_47),.clk(clk),.wout(w18_47));
	PE pe18_48(.x(x48),.w(w18_47),.acc(r18_47),.res(r18_48),.clk(clk),.wout(w18_48));
	PE pe18_49(.x(x49),.w(w18_48),.acc(r18_48),.res(r18_49),.clk(clk),.wout(w18_49));
	PE pe18_50(.x(x50),.w(w18_49),.acc(r18_49),.res(r18_50),.clk(clk),.wout(w18_50));
	PE pe18_51(.x(x51),.w(w18_50),.acc(r18_50),.res(r18_51),.clk(clk),.wout(w18_51));
	PE pe18_52(.x(x52),.w(w18_51),.acc(r18_51),.res(r18_52),.clk(clk),.wout(w18_52));
	PE pe18_53(.x(x53),.w(w18_52),.acc(r18_52),.res(r18_53),.clk(clk),.wout(w18_53));
	PE pe18_54(.x(x54),.w(w18_53),.acc(r18_53),.res(r18_54),.clk(clk),.wout(w18_54));
	PE pe18_55(.x(x55),.w(w18_54),.acc(r18_54),.res(r18_55),.clk(clk),.wout(w18_55));
	PE pe18_56(.x(x56),.w(w18_55),.acc(r18_55),.res(r18_56),.clk(clk),.wout(w18_56));
	PE pe18_57(.x(x57),.w(w18_56),.acc(r18_56),.res(r18_57),.clk(clk),.wout(w18_57));
	PE pe18_58(.x(x58),.w(w18_57),.acc(r18_57),.res(r18_58),.clk(clk),.wout(w18_58));
	PE pe18_59(.x(x59),.w(w18_58),.acc(r18_58),.res(r18_59),.clk(clk),.wout(w18_59));
	PE pe18_60(.x(x60),.w(w18_59),.acc(r18_59),.res(r18_60),.clk(clk),.wout(w18_60));
	PE pe18_61(.x(x61),.w(w18_60),.acc(r18_60),.res(r18_61),.clk(clk),.wout(w18_61));
	PE pe18_62(.x(x62),.w(w18_61),.acc(r18_61),.res(r18_62),.clk(clk),.wout(w18_62));
	PE pe18_63(.x(x63),.w(w18_62),.acc(r18_62),.res(r18_63),.clk(clk),.wout(w18_63));
	PE pe18_64(.x(x64),.w(w18_63),.acc(r18_63),.res(r18_64),.clk(clk),.wout(w18_64));
	PE pe18_65(.x(x65),.w(w18_64),.acc(r18_64),.res(r18_65),.clk(clk),.wout(w18_65));
	PE pe18_66(.x(x66),.w(w18_65),.acc(r18_65),.res(r18_66),.clk(clk),.wout(w18_66));
	PE pe18_67(.x(x67),.w(w18_66),.acc(r18_66),.res(r18_67),.clk(clk),.wout(w18_67));
	PE pe18_68(.x(x68),.w(w18_67),.acc(r18_67),.res(r18_68),.clk(clk),.wout(w18_68));
	PE pe18_69(.x(x69),.w(w18_68),.acc(r18_68),.res(r18_69),.clk(clk),.wout(w18_69));
	PE pe18_70(.x(x70),.w(w18_69),.acc(r18_69),.res(r18_70),.clk(clk),.wout(w18_70));
	PE pe18_71(.x(x71),.w(w18_70),.acc(r18_70),.res(r18_71),.clk(clk),.wout(w18_71));
	PE pe18_72(.x(x72),.w(w18_71),.acc(r18_71),.res(r18_72),.clk(clk),.wout(w18_72));
	PE pe18_73(.x(x73),.w(w18_72),.acc(r18_72),.res(r18_73),.clk(clk),.wout(w18_73));
	PE pe18_74(.x(x74),.w(w18_73),.acc(r18_73),.res(r18_74),.clk(clk),.wout(w18_74));
	PE pe18_75(.x(x75),.w(w18_74),.acc(r18_74),.res(r18_75),.clk(clk),.wout(w18_75));
	PE pe18_76(.x(x76),.w(w18_75),.acc(r18_75),.res(r18_76),.clk(clk),.wout(w18_76));
	PE pe18_77(.x(x77),.w(w18_76),.acc(r18_76),.res(r18_77),.clk(clk),.wout(w18_77));
	PE pe18_78(.x(x78),.w(w18_77),.acc(r18_77),.res(r18_78),.clk(clk),.wout(w18_78));
	PE pe18_79(.x(x79),.w(w18_78),.acc(r18_78),.res(r18_79),.clk(clk),.wout(w18_79));
	PE pe18_80(.x(x80),.w(w18_79),.acc(r18_79),.res(r18_80),.clk(clk),.wout(w18_80));
	PE pe18_81(.x(x81),.w(w18_80),.acc(r18_80),.res(r18_81),.clk(clk),.wout(w18_81));
	PE pe18_82(.x(x82),.w(w18_81),.acc(r18_81),.res(r18_82),.clk(clk),.wout(w18_82));
	PE pe18_83(.x(x83),.w(w18_82),.acc(r18_82),.res(r18_83),.clk(clk),.wout(w18_83));
	PE pe18_84(.x(x84),.w(w18_83),.acc(r18_83),.res(r18_84),.clk(clk),.wout(w18_84));
	PE pe18_85(.x(x85),.w(w18_84),.acc(r18_84),.res(r18_85),.clk(clk),.wout(w18_85));
	PE pe18_86(.x(x86),.w(w18_85),.acc(r18_85),.res(r18_86),.clk(clk),.wout(w18_86));
	PE pe18_87(.x(x87),.w(w18_86),.acc(r18_86),.res(r18_87),.clk(clk),.wout(w18_87));
	PE pe18_88(.x(x88),.w(w18_87),.acc(r18_87),.res(r18_88),.clk(clk),.wout(w18_88));
	PE pe18_89(.x(x89),.w(w18_88),.acc(r18_88),.res(r18_89),.clk(clk),.wout(w18_89));
	PE pe18_90(.x(x90),.w(w18_89),.acc(r18_89),.res(r18_90),.clk(clk),.wout(w18_90));
	PE pe18_91(.x(x91),.w(w18_90),.acc(r18_90),.res(r18_91),.clk(clk),.wout(w18_91));
	PE pe18_92(.x(x92),.w(w18_91),.acc(r18_91),.res(r18_92),.clk(clk),.wout(w18_92));
	PE pe18_93(.x(x93),.w(w18_92),.acc(r18_92),.res(r18_93),.clk(clk),.wout(w18_93));
	PE pe18_94(.x(x94),.w(w18_93),.acc(r18_93),.res(r18_94),.clk(clk),.wout(w18_94));
	PE pe18_95(.x(x95),.w(w18_94),.acc(r18_94),.res(r18_95),.clk(clk),.wout(w18_95));
	PE pe18_96(.x(x96),.w(w18_95),.acc(r18_95),.res(r18_96),.clk(clk),.wout(w18_96));
	PE pe18_97(.x(x97),.w(w18_96),.acc(r18_96),.res(r18_97),.clk(clk),.wout(w18_97));
	PE pe18_98(.x(x98),.w(w18_97),.acc(r18_97),.res(r18_98),.clk(clk),.wout(w18_98));
	PE pe18_99(.x(x99),.w(w18_98),.acc(r18_98),.res(r18_99),.clk(clk),.wout(w18_99));
	PE pe18_100(.x(x100),.w(w18_99),.acc(r18_99),.res(r18_100),.clk(clk),.wout(w18_100));
	PE pe18_101(.x(x101),.w(w18_100),.acc(r18_100),.res(r18_101),.clk(clk),.wout(w18_101));
	PE pe18_102(.x(x102),.w(w18_101),.acc(r18_101),.res(r18_102),.clk(clk),.wout(w18_102));
	PE pe18_103(.x(x103),.w(w18_102),.acc(r18_102),.res(r18_103),.clk(clk),.wout(w18_103));
	PE pe18_104(.x(x104),.w(w18_103),.acc(r18_103),.res(r18_104),.clk(clk),.wout(w18_104));
	PE pe18_105(.x(x105),.w(w18_104),.acc(r18_104),.res(r18_105),.clk(clk),.wout(w18_105));
	PE pe18_106(.x(x106),.w(w18_105),.acc(r18_105),.res(r18_106),.clk(clk),.wout(w18_106));
	PE pe18_107(.x(x107),.w(w18_106),.acc(r18_106),.res(r18_107),.clk(clk),.wout(w18_107));
	PE pe18_108(.x(x108),.w(w18_107),.acc(r18_107),.res(r18_108),.clk(clk),.wout(w18_108));
	PE pe18_109(.x(x109),.w(w18_108),.acc(r18_108),.res(r18_109),.clk(clk),.wout(w18_109));
	PE pe18_110(.x(x110),.w(w18_109),.acc(r18_109),.res(r18_110),.clk(clk),.wout(w18_110));
	PE pe18_111(.x(x111),.w(w18_110),.acc(r18_110),.res(r18_111),.clk(clk),.wout(w18_111));
	PE pe18_112(.x(x112),.w(w18_111),.acc(r18_111),.res(r18_112),.clk(clk),.wout(w18_112));
	PE pe18_113(.x(x113),.w(w18_112),.acc(r18_112),.res(r18_113),.clk(clk),.wout(w18_113));
	PE pe18_114(.x(x114),.w(w18_113),.acc(r18_113),.res(r18_114),.clk(clk),.wout(w18_114));
	PE pe18_115(.x(x115),.w(w18_114),.acc(r18_114),.res(r18_115),.clk(clk),.wout(w18_115));
	PE pe18_116(.x(x116),.w(w18_115),.acc(r18_115),.res(r18_116),.clk(clk),.wout(w18_116));
	PE pe18_117(.x(x117),.w(w18_116),.acc(r18_116),.res(r18_117),.clk(clk),.wout(w18_117));
	PE pe18_118(.x(x118),.w(w18_117),.acc(r18_117),.res(r18_118),.clk(clk),.wout(w18_118));
	PE pe18_119(.x(x119),.w(w18_118),.acc(r18_118),.res(r18_119),.clk(clk),.wout(w18_119));
	PE pe18_120(.x(x120),.w(w18_119),.acc(r18_119),.res(r18_120),.clk(clk),.wout(w18_120));
	PE pe18_121(.x(x121),.w(w18_120),.acc(r18_120),.res(r18_121),.clk(clk),.wout(w18_121));
	PE pe18_122(.x(x122),.w(w18_121),.acc(r18_121),.res(r18_122),.clk(clk),.wout(w18_122));
	PE pe18_123(.x(x123),.w(w18_122),.acc(r18_122),.res(r18_123),.clk(clk),.wout(w18_123));
	PE pe18_124(.x(x124),.w(w18_123),.acc(r18_123),.res(r18_124),.clk(clk),.wout(w18_124));
	PE pe18_125(.x(x125),.w(w18_124),.acc(r18_124),.res(r18_125),.clk(clk),.wout(w18_125));
	PE pe18_126(.x(x126),.w(w18_125),.acc(r18_125),.res(r18_126),.clk(clk),.wout(w18_126));
	PE pe18_127(.x(x127),.w(w18_126),.acc(r18_126),.res(result18),.clk(clk),.wout(weight18));

	PE pe19_0(.x(x0),.w(w19),.acc(32'h0),.res(r19_0),.clk(clk),.wout(w19_0));
	PE pe19_1(.x(x1),.w(w19_0),.acc(r19_0),.res(r19_1),.clk(clk),.wout(w19_1));
	PE pe19_2(.x(x2),.w(w19_1),.acc(r19_1),.res(r19_2),.clk(clk),.wout(w19_2));
	PE pe19_3(.x(x3),.w(w19_2),.acc(r19_2),.res(r19_3),.clk(clk),.wout(w19_3));
	PE pe19_4(.x(x4),.w(w19_3),.acc(r19_3),.res(r19_4),.clk(clk),.wout(w19_4));
	PE pe19_5(.x(x5),.w(w19_4),.acc(r19_4),.res(r19_5),.clk(clk),.wout(w19_5));
	PE pe19_6(.x(x6),.w(w19_5),.acc(r19_5),.res(r19_6),.clk(clk),.wout(w19_6));
	PE pe19_7(.x(x7),.w(w19_6),.acc(r19_6),.res(r19_7),.clk(clk),.wout(w19_7));
	PE pe19_8(.x(x8),.w(w19_7),.acc(r19_7),.res(r19_8),.clk(clk),.wout(w19_8));
	PE pe19_9(.x(x9),.w(w19_8),.acc(r19_8),.res(r19_9),.clk(clk),.wout(w19_9));
	PE pe19_10(.x(x10),.w(w19_9),.acc(r19_9),.res(r19_10),.clk(clk),.wout(w19_10));
	PE pe19_11(.x(x11),.w(w19_10),.acc(r19_10),.res(r19_11),.clk(clk),.wout(w19_11));
	PE pe19_12(.x(x12),.w(w19_11),.acc(r19_11),.res(r19_12),.clk(clk),.wout(w19_12));
	PE pe19_13(.x(x13),.w(w19_12),.acc(r19_12),.res(r19_13),.clk(clk),.wout(w19_13));
	PE pe19_14(.x(x14),.w(w19_13),.acc(r19_13),.res(r19_14),.clk(clk),.wout(w19_14));
	PE pe19_15(.x(x15),.w(w19_14),.acc(r19_14),.res(r19_15),.clk(clk),.wout(w19_15));
	PE pe19_16(.x(x16),.w(w19_15),.acc(r19_15),.res(r19_16),.clk(clk),.wout(w19_16));
	PE pe19_17(.x(x17),.w(w19_16),.acc(r19_16),.res(r19_17),.clk(clk),.wout(w19_17));
	PE pe19_18(.x(x18),.w(w19_17),.acc(r19_17),.res(r19_18),.clk(clk),.wout(w19_18));
	PE pe19_19(.x(x19),.w(w19_18),.acc(r19_18),.res(r19_19),.clk(clk),.wout(w19_19));
	PE pe19_20(.x(x20),.w(w19_19),.acc(r19_19),.res(r19_20),.clk(clk),.wout(w19_20));
	PE pe19_21(.x(x21),.w(w19_20),.acc(r19_20),.res(r19_21),.clk(clk),.wout(w19_21));
	PE pe19_22(.x(x22),.w(w19_21),.acc(r19_21),.res(r19_22),.clk(clk),.wout(w19_22));
	PE pe19_23(.x(x23),.w(w19_22),.acc(r19_22),.res(r19_23),.clk(clk),.wout(w19_23));
	PE pe19_24(.x(x24),.w(w19_23),.acc(r19_23),.res(r19_24),.clk(clk),.wout(w19_24));
	PE pe19_25(.x(x25),.w(w19_24),.acc(r19_24),.res(r19_25),.clk(clk),.wout(w19_25));
	PE pe19_26(.x(x26),.w(w19_25),.acc(r19_25),.res(r19_26),.clk(clk),.wout(w19_26));
	PE pe19_27(.x(x27),.w(w19_26),.acc(r19_26),.res(r19_27),.clk(clk),.wout(w19_27));
	PE pe19_28(.x(x28),.w(w19_27),.acc(r19_27),.res(r19_28),.clk(clk),.wout(w19_28));
	PE pe19_29(.x(x29),.w(w19_28),.acc(r19_28),.res(r19_29),.clk(clk),.wout(w19_29));
	PE pe19_30(.x(x30),.w(w19_29),.acc(r19_29),.res(r19_30),.clk(clk),.wout(w19_30));
	PE pe19_31(.x(x31),.w(w19_30),.acc(r19_30),.res(r19_31),.clk(clk),.wout(w19_31));
	PE pe19_32(.x(x32),.w(w19_31),.acc(r19_31),.res(r19_32),.clk(clk),.wout(w19_32));
	PE pe19_33(.x(x33),.w(w19_32),.acc(r19_32),.res(r19_33),.clk(clk),.wout(w19_33));
	PE pe19_34(.x(x34),.w(w19_33),.acc(r19_33),.res(r19_34),.clk(clk),.wout(w19_34));
	PE pe19_35(.x(x35),.w(w19_34),.acc(r19_34),.res(r19_35),.clk(clk),.wout(w19_35));
	PE pe19_36(.x(x36),.w(w19_35),.acc(r19_35),.res(r19_36),.clk(clk),.wout(w19_36));
	PE pe19_37(.x(x37),.w(w19_36),.acc(r19_36),.res(r19_37),.clk(clk),.wout(w19_37));
	PE pe19_38(.x(x38),.w(w19_37),.acc(r19_37),.res(r19_38),.clk(clk),.wout(w19_38));
	PE pe19_39(.x(x39),.w(w19_38),.acc(r19_38),.res(r19_39),.clk(clk),.wout(w19_39));
	PE pe19_40(.x(x40),.w(w19_39),.acc(r19_39),.res(r19_40),.clk(clk),.wout(w19_40));
	PE pe19_41(.x(x41),.w(w19_40),.acc(r19_40),.res(r19_41),.clk(clk),.wout(w19_41));
	PE pe19_42(.x(x42),.w(w19_41),.acc(r19_41),.res(r19_42),.clk(clk),.wout(w19_42));
	PE pe19_43(.x(x43),.w(w19_42),.acc(r19_42),.res(r19_43),.clk(clk),.wout(w19_43));
	PE pe19_44(.x(x44),.w(w19_43),.acc(r19_43),.res(r19_44),.clk(clk),.wout(w19_44));
	PE pe19_45(.x(x45),.w(w19_44),.acc(r19_44),.res(r19_45),.clk(clk),.wout(w19_45));
	PE pe19_46(.x(x46),.w(w19_45),.acc(r19_45),.res(r19_46),.clk(clk),.wout(w19_46));
	PE pe19_47(.x(x47),.w(w19_46),.acc(r19_46),.res(r19_47),.clk(clk),.wout(w19_47));
	PE pe19_48(.x(x48),.w(w19_47),.acc(r19_47),.res(r19_48),.clk(clk),.wout(w19_48));
	PE pe19_49(.x(x49),.w(w19_48),.acc(r19_48),.res(r19_49),.clk(clk),.wout(w19_49));
	PE pe19_50(.x(x50),.w(w19_49),.acc(r19_49),.res(r19_50),.clk(clk),.wout(w19_50));
	PE pe19_51(.x(x51),.w(w19_50),.acc(r19_50),.res(r19_51),.clk(clk),.wout(w19_51));
	PE pe19_52(.x(x52),.w(w19_51),.acc(r19_51),.res(r19_52),.clk(clk),.wout(w19_52));
	PE pe19_53(.x(x53),.w(w19_52),.acc(r19_52),.res(r19_53),.clk(clk),.wout(w19_53));
	PE pe19_54(.x(x54),.w(w19_53),.acc(r19_53),.res(r19_54),.clk(clk),.wout(w19_54));
	PE pe19_55(.x(x55),.w(w19_54),.acc(r19_54),.res(r19_55),.clk(clk),.wout(w19_55));
	PE pe19_56(.x(x56),.w(w19_55),.acc(r19_55),.res(r19_56),.clk(clk),.wout(w19_56));
	PE pe19_57(.x(x57),.w(w19_56),.acc(r19_56),.res(r19_57),.clk(clk),.wout(w19_57));
	PE pe19_58(.x(x58),.w(w19_57),.acc(r19_57),.res(r19_58),.clk(clk),.wout(w19_58));
	PE pe19_59(.x(x59),.w(w19_58),.acc(r19_58),.res(r19_59),.clk(clk),.wout(w19_59));
	PE pe19_60(.x(x60),.w(w19_59),.acc(r19_59),.res(r19_60),.clk(clk),.wout(w19_60));
	PE pe19_61(.x(x61),.w(w19_60),.acc(r19_60),.res(r19_61),.clk(clk),.wout(w19_61));
	PE pe19_62(.x(x62),.w(w19_61),.acc(r19_61),.res(r19_62),.clk(clk),.wout(w19_62));
	PE pe19_63(.x(x63),.w(w19_62),.acc(r19_62),.res(r19_63),.clk(clk),.wout(w19_63));
	PE pe19_64(.x(x64),.w(w19_63),.acc(r19_63),.res(r19_64),.clk(clk),.wout(w19_64));
	PE pe19_65(.x(x65),.w(w19_64),.acc(r19_64),.res(r19_65),.clk(clk),.wout(w19_65));
	PE pe19_66(.x(x66),.w(w19_65),.acc(r19_65),.res(r19_66),.clk(clk),.wout(w19_66));
	PE pe19_67(.x(x67),.w(w19_66),.acc(r19_66),.res(r19_67),.clk(clk),.wout(w19_67));
	PE pe19_68(.x(x68),.w(w19_67),.acc(r19_67),.res(r19_68),.clk(clk),.wout(w19_68));
	PE pe19_69(.x(x69),.w(w19_68),.acc(r19_68),.res(r19_69),.clk(clk),.wout(w19_69));
	PE pe19_70(.x(x70),.w(w19_69),.acc(r19_69),.res(r19_70),.clk(clk),.wout(w19_70));
	PE pe19_71(.x(x71),.w(w19_70),.acc(r19_70),.res(r19_71),.clk(clk),.wout(w19_71));
	PE pe19_72(.x(x72),.w(w19_71),.acc(r19_71),.res(r19_72),.clk(clk),.wout(w19_72));
	PE pe19_73(.x(x73),.w(w19_72),.acc(r19_72),.res(r19_73),.clk(clk),.wout(w19_73));
	PE pe19_74(.x(x74),.w(w19_73),.acc(r19_73),.res(r19_74),.clk(clk),.wout(w19_74));
	PE pe19_75(.x(x75),.w(w19_74),.acc(r19_74),.res(r19_75),.clk(clk),.wout(w19_75));
	PE pe19_76(.x(x76),.w(w19_75),.acc(r19_75),.res(r19_76),.clk(clk),.wout(w19_76));
	PE pe19_77(.x(x77),.w(w19_76),.acc(r19_76),.res(r19_77),.clk(clk),.wout(w19_77));
	PE pe19_78(.x(x78),.w(w19_77),.acc(r19_77),.res(r19_78),.clk(clk),.wout(w19_78));
	PE pe19_79(.x(x79),.w(w19_78),.acc(r19_78),.res(r19_79),.clk(clk),.wout(w19_79));
	PE pe19_80(.x(x80),.w(w19_79),.acc(r19_79),.res(r19_80),.clk(clk),.wout(w19_80));
	PE pe19_81(.x(x81),.w(w19_80),.acc(r19_80),.res(r19_81),.clk(clk),.wout(w19_81));
	PE pe19_82(.x(x82),.w(w19_81),.acc(r19_81),.res(r19_82),.clk(clk),.wout(w19_82));
	PE pe19_83(.x(x83),.w(w19_82),.acc(r19_82),.res(r19_83),.clk(clk),.wout(w19_83));
	PE pe19_84(.x(x84),.w(w19_83),.acc(r19_83),.res(r19_84),.clk(clk),.wout(w19_84));
	PE pe19_85(.x(x85),.w(w19_84),.acc(r19_84),.res(r19_85),.clk(clk),.wout(w19_85));
	PE pe19_86(.x(x86),.w(w19_85),.acc(r19_85),.res(r19_86),.clk(clk),.wout(w19_86));
	PE pe19_87(.x(x87),.w(w19_86),.acc(r19_86),.res(r19_87),.clk(clk),.wout(w19_87));
	PE pe19_88(.x(x88),.w(w19_87),.acc(r19_87),.res(r19_88),.clk(clk),.wout(w19_88));
	PE pe19_89(.x(x89),.w(w19_88),.acc(r19_88),.res(r19_89),.clk(clk),.wout(w19_89));
	PE pe19_90(.x(x90),.w(w19_89),.acc(r19_89),.res(r19_90),.clk(clk),.wout(w19_90));
	PE pe19_91(.x(x91),.w(w19_90),.acc(r19_90),.res(r19_91),.clk(clk),.wout(w19_91));
	PE pe19_92(.x(x92),.w(w19_91),.acc(r19_91),.res(r19_92),.clk(clk),.wout(w19_92));
	PE pe19_93(.x(x93),.w(w19_92),.acc(r19_92),.res(r19_93),.clk(clk),.wout(w19_93));
	PE pe19_94(.x(x94),.w(w19_93),.acc(r19_93),.res(r19_94),.clk(clk),.wout(w19_94));
	PE pe19_95(.x(x95),.w(w19_94),.acc(r19_94),.res(r19_95),.clk(clk),.wout(w19_95));
	PE pe19_96(.x(x96),.w(w19_95),.acc(r19_95),.res(r19_96),.clk(clk),.wout(w19_96));
	PE pe19_97(.x(x97),.w(w19_96),.acc(r19_96),.res(r19_97),.clk(clk),.wout(w19_97));
	PE pe19_98(.x(x98),.w(w19_97),.acc(r19_97),.res(r19_98),.clk(clk),.wout(w19_98));
	PE pe19_99(.x(x99),.w(w19_98),.acc(r19_98),.res(r19_99),.clk(clk),.wout(w19_99));
	PE pe19_100(.x(x100),.w(w19_99),.acc(r19_99),.res(r19_100),.clk(clk),.wout(w19_100));
	PE pe19_101(.x(x101),.w(w19_100),.acc(r19_100),.res(r19_101),.clk(clk),.wout(w19_101));
	PE pe19_102(.x(x102),.w(w19_101),.acc(r19_101),.res(r19_102),.clk(clk),.wout(w19_102));
	PE pe19_103(.x(x103),.w(w19_102),.acc(r19_102),.res(r19_103),.clk(clk),.wout(w19_103));
	PE pe19_104(.x(x104),.w(w19_103),.acc(r19_103),.res(r19_104),.clk(clk),.wout(w19_104));
	PE pe19_105(.x(x105),.w(w19_104),.acc(r19_104),.res(r19_105),.clk(clk),.wout(w19_105));
	PE pe19_106(.x(x106),.w(w19_105),.acc(r19_105),.res(r19_106),.clk(clk),.wout(w19_106));
	PE pe19_107(.x(x107),.w(w19_106),.acc(r19_106),.res(r19_107),.clk(clk),.wout(w19_107));
	PE pe19_108(.x(x108),.w(w19_107),.acc(r19_107),.res(r19_108),.clk(clk),.wout(w19_108));
	PE pe19_109(.x(x109),.w(w19_108),.acc(r19_108),.res(r19_109),.clk(clk),.wout(w19_109));
	PE pe19_110(.x(x110),.w(w19_109),.acc(r19_109),.res(r19_110),.clk(clk),.wout(w19_110));
	PE pe19_111(.x(x111),.w(w19_110),.acc(r19_110),.res(r19_111),.clk(clk),.wout(w19_111));
	PE pe19_112(.x(x112),.w(w19_111),.acc(r19_111),.res(r19_112),.clk(clk),.wout(w19_112));
	PE pe19_113(.x(x113),.w(w19_112),.acc(r19_112),.res(r19_113),.clk(clk),.wout(w19_113));
	PE pe19_114(.x(x114),.w(w19_113),.acc(r19_113),.res(r19_114),.clk(clk),.wout(w19_114));
	PE pe19_115(.x(x115),.w(w19_114),.acc(r19_114),.res(r19_115),.clk(clk),.wout(w19_115));
	PE pe19_116(.x(x116),.w(w19_115),.acc(r19_115),.res(r19_116),.clk(clk),.wout(w19_116));
	PE pe19_117(.x(x117),.w(w19_116),.acc(r19_116),.res(r19_117),.clk(clk),.wout(w19_117));
	PE pe19_118(.x(x118),.w(w19_117),.acc(r19_117),.res(r19_118),.clk(clk),.wout(w19_118));
	PE pe19_119(.x(x119),.w(w19_118),.acc(r19_118),.res(r19_119),.clk(clk),.wout(w19_119));
	PE pe19_120(.x(x120),.w(w19_119),.acc(r19_119),.res(r19_120),.clk(clk),.wout(w19_120));
	PE pe19_121(.x(x121),.w(w19_120),.acc(r19_120),.res(r19_121),.clk(clk),.wout(w19_121));
	PE pe19_122(.x(x122),.w(w19_121),.acc(r19_121),.res(r19_122),.clk(clk),.wout(w19_122));
	PE pe19_123(.x(x123),.w(w19_122),.acc(r19_122),.res(r19_123),.clk(clk),.wout(w19_123));
	PE pe19_124(.x(x124),.w(w19_123),.acc(r19_123),.res(r19_124),.clk(clk),.wout(w19_124));
	PE pe19_125(.x(x125),.w(w19_124),.acc(r19_124),.res(r19_125),.clk(clk),.wout(w19_125));
	PE pe19_126(.x(x126),.w(w19_125),.acc(r19_125),.res(r19_126),.clk(clk),.wout(w19_126));
	PE pe19_127(.x(x127),.w(w19_126),.acc(r19_126),.res(result19),.clk(clk),.wout(weight19));

	PE pe20_0(.x(x0),.w(w20),.acc(32'h0),.res(r20_0),.clk(clk),.wout(w20_0));
	PE pe20_1(.x(x1),.w(w20_0),.acc(r20_0),.res(r20_1),.clk(clk),.wout(w20_1));
	PE pe20_2(.x(x2),.w(w20_1),.acc(r20_1),.res(r20_2),.clk(clk),.wout(w20_2));
	PE pe20_3(.x(x3),.w(w20_2),.acc(r20_2),.res(r20_3),.clk(clk),.wout(w20_3));
	PE pe20_4(.x(x4),.w(w20_3),.acc(r20_3),.res(r20_4),.clk(clk),.wout(w20_4));
	PE pe20_5(.x(x5),.w(w20_4),.acc(r20_4),.res(r20_5),.clk(clk),.wout(w20_5));
	PE pe20_6(.x(x6),.w(w20_5),.acc(r20_5),.res(r20_6),.clk(clk),.wout(w20_6));
	PE pe20_7(.x(x7),.w(w20_6),.acc(r20_6),.res(r20_7),.clk(clk),.wout(w20_7));
	PE pe20_8(.x(x8),.w(w20_7),.acc(r20_7),.res(r20_8),.clk(clk),.wout(w20_8));
	PE pe20_9(.x(x9),.w(w20_8),.acc(r20_8),.res(r20_9),.clk(clk),.wout(w20_9));
	PE pe20_10(.x(x10),.w(w20_9),.acc(r20_9),.res(r20_10),.clk(clk),.wout(w20_10));
	PE pe20_11(.x(x11),.w(w20_10),.acc(r20_10),.res(r20_11),.clk(clk),.wout(w20_11));
	PE pe20_12(.x(x12),.w(w20_11),.acc(r20_11),.res(r20_12),.clk(clk),.wout(w20_12));
	PE pe20_13(.x(x13),.w(w20_12),.acc(r20_12),.res(r20_13),.clk(clk),.wout(w20_13));
	PE pe20_14(.x(x14),.w(w20_13),.acc(r20_13),.res(r20_14),.clk(clk),.wout(w20_14));
	PE pe20_15(.x(x15),.w(w20_14),.acc(r20_14),.res(r20_15),.clk(clk),.wout(w20_15));
	PE pe20_16(.x(x16),.w(w20_15),.acc(r20_15),.res(r20_16),.clk(clk),.wout(w20_16));
	PE pe20_17(.x(x17),.w(w20_16),.acc(r20_16),.res(r20_17),.clk(clk),.wout(w20_17));
	PE pe20_18(.x(x18),.w(w20_17),.acc(r20_17),.res(r20_18),.clk(clk),.wout(w20_18));
	PE pe20_19(.x(x19),.w(w20_18),.acc(r20_18),.res(r20_19),.clk(clk),.wout(w20_19));
	PE pe20_20(.x(x20),.w(w20_19),.acc(r20_19),.res(r20_20),.clk(clk),.wout(w20_20));
	PE pe20_21(.x(x21),.w(w20_20),.acc(r20_20),.res(r20_21),.clk(clk),.wout(w20_21));
	PE pe20_22(.x(x22),.w(w20_21),.acc(r20_21),.res(r20_22),.clk(clk),.wout(w20_22));
	PE pe20_23(.x(x23),.w(w20_22),.acc(r20_22),.res(r20_23),.clk(clk),.wout(w20_23));
	PE pe20_24(.x(x24),.w(w20_23),.acc(r20_23),.res(r20_24),.clk(clk),.wout(w20_24));
	PE pe20_25(.x(x25),.w(w20_24),.acc(r20_24),.res(r20_25),.clk(clk),.wout(w20_25));
	PE pe20_26(.x(x26),.w(w20_25),.acc(r20_25),.res(r20_26),.clk(clk),.wout(w20_26));
	PE pe20_27(.x(x27),.w(w20_26),.acc(r20_26),.res(r20_27),.clk(clk),.wout(w20_27));
	PE pe20_28(.x(x28),.w(w20_27),.acc(r20_27),.res(r20_28),.clk(clk),.wout(w20_28));
	PE pe20_29(.x(x29),.w(w20_28),.acc(r20_28),.res(r20_29),.clk(clk),.wout(w20_29));
	PE pe20_30(.x(x30),.w(w20_29),.acc(r20_29),.res(r20_30),.clk(clk),.wout(w20_30));
	PE pe20_31(.x(x31),.w(w20_30),.acc(r20_30),.res(r20_31),.clk(clk),.wout(w20_31));
	PE pe20_32(.x(x32),.w(w20_31),.acc(r20_31),.res(r20_32),.clk(clk),.wout(w20_32));
	PE pe20_33(.x(x33),.w(w20_32),.acc(r20_32),.res(r20_33),.clk(clk),.wout(w20_33));
	PE pe20_34(.x(x34),.w(w20_33),.acc(r20_33),.res(r20_34),.clk(clk),.wout(w20_34));
	PE pe20_35(.x(x35),.w(w20_34),.acc(r20_34),.res(r20_35),.clk(clk),.wout(w20_35));
	PE pe20_36(.x(x36),.w(w20_35),.acc(r20_35),.res(r20_36),.clk(clk),.wout(w20_36));
	PE pe20_37(.x(x37),.w(w20_36),.acc(r20_36),.res(r20_37),.clk(clk),.wout(w20_37));
	PE pe20_38(.x(x38),.w(w20_37),.acc(r20_37),.res(r20_38),.clk(clk),.wout(w20_38));
	PE pe20_39(.x(x39),.w(w20_38),.acc(r20_38),.res(r20_39),.clk(clk),.wout(w20_39));
	PE pe20_40(.x(x40),.w(w20_39),.acc(r20_39),.res(r20_40),.clk(clk),.wout(w20_40));
	PE pe20_41(.x(x41),.w(w20_40),.acc(r20_40),.res(r20_41),.clk(clk),.wout(w20_41));
	PE pe20_42(.x(x42),.w(w20_41),.acc(r20_41),.res(r20_42),.clk(clk),.wout(w20_42));
	PE pe20_43(.x(x43),.w(w20_42),.acc(r20_42),.res(r20_43),.clk(clk),.wout(w20_43));
	PE pe20_44(.x(x44),.w(w20_43),.acc(r20_43),.res(r20_44),.clk(clk),.wout(w20_44));
	PE pe20_45(.x(x45),.w(w20_44),.acc(r20_44),.res(r20_45),.clk(clk),.wout(w20_45));
	PE pe20_46(.x(x46),.w(w20_45),.acc(r20_45),.res(r20_46),.clk(clk),.wout(w20_46));
	PE pe20_47(.x(x47),.w(w20_46),.acc(r20_46),.res(r20_47),.clk(clk),.wout(w20_47));
	PE pe20_48(.x(x48),.w(w20_47),.acc(r20_47),.res(r20_48),.clk(clk),.wout(w20_48));
	PE pe20_49(.x(x49),.w(w20_48),.acc(r20_48),.res(r20_49),.clk(clk),.wout(w20_49));
	PE pe20_50(.x(x50),.w(w20_49),.acc(r20_49),.res(r20_50),.clk(clk),.wout(w20_50));
	PE pe20_51(.x(x51),.w(w20_50),.acc(r20_50),.res(r20_51),.clk(clk),.wout(w20_51));
	PE pe20_52(.x(x52),.w(w20_51),.acc(r20_51),.res(r20_52),.clk(clk),.wout(w20_52));
	PE pe20_53(.x(x53),.w(w20_52),.acc(r20_52),.res(r20_53),.clk(clk),.wout(w20_53));
	PE pe20_54(.x(x54),.w(w20_53),.acc(r20_53),.res(r20_54),.clk(clk),.wout(w20_54));
	PE pe20_55(.x(x55),.w(w20_54),.acc(r20_54),.res(r20_55),.clk(clk),.wout(w20_55));
	PE pe20_56(.x(x56),.w(w20_55),.acc(r20_55),.res(r20_56),.clk(clk),.wout(w20_56));
	PE pe20_57(.x(x57),.w(w20_56),.acc(r20_56),.res(r20_57),.clk(clk),.wout(w20_57));
	PE pe20_58(.x(x58),.w(w20_57),.acc(r20_57),.res(r20_58),.clk(clk),.wout(w20_58));
	PE pe20_59(.x(x59),.w(w20_58),.acc(r20_58),.res(r20_59),.clk(clk),.wout(w20_59));
	PE pe20_60(.x(x60),.w(w20_59),.acc(r20_59),.res(r20_60),.clk(clk),.wout(w20_60));
	PE pe20_61(.x(x61),.w(w20_60),.acc(r20_60),.res(r20_61),.clk(clk),.wout(w20_61));
	PE pe20_62(.x(x62),.w(w20_61),.acc(r20_61),.res(r20_62),.clk(clk),.wout(w20_62));
	PE pe20_63(.x(x63),.w(w20_62),.acc(r20_62),.res(r20_63),.clk(clk),.wout(w20_63));
	PE pe20_64(.x(x64),.w(w20_63),.acc(r20_63),.res(r20_64),.clk(clk),.wout(w20_64));
	PE pe20_65(.x(x65),.w(w20_64),.acc(r20_64),.res(r20_65),.clk(clk),.wout(w20_65));
	PE pe20_66(.x(x66),.w(w20_65),.acc(r20_65),.res(r20_66),.clk(clk),.wout(w20_66));
	PE pe20_67(.x(x67),.w(w20_66),.acc(r20_66),.res(r20_67),.clk(clk),.wout(w20_67));
	PE pe20_68(.x(x68),.w(w20_67),.acc(r20_67),.res(r20_68),.clk(clk),.wout(w20_68));
	PE pe20_69(.x(x69),.w(w20_68),.acc(r20_68),.res(r20_69),.clk(clk),.wout(w20_69));
	PE pe20_70(.x(x70),.w(w20_69),.acc(r20_69),.res(r20_70),.clk(clk),.wout(w20_70));
	PE pe20_71(.x(x71),.w(w20_70),.acc(r20_70),.res(r20_71),.clk(clk),.wout(w20_71));
	PE pe20_72(.x(x72),.w(w20_71),.acc(r20_71),.res(r20_72),.clk(clk),.wout(w20_72));
	PE pe20_73(.x(x73),.w(w20_72),.acc(r20_72),.res(r20_73),.clk(clk),.wout(w20_73));
	PE pe20_74(.x(x74),.w(w20_73),.acc(r20_73),.res(r20_74),.clk(clk),.wout(w20_74));
	PE pe20_75(.x(x75),.w(w20_74),.acc(r20_74),.res(r20_75),.clk(clk),.wout(w20_75));
	PE pe20_76(.x(x76),.w(w20_75),.acc(r20_75),.res(r20_76),.clk(clk),.wout(w20_76));
	PE pe20_77(.x(x77),.w(w20_76),.acc(r20_76),.res(r20_77),.clk(clk),.wout(w20_77));
	PE pe20_78(.x(x78),.w(w20_77),.acc(r20_77),.res(r20_78),.clk(clk),.wout(w20_78));
	PE pe20_79(.x(x79),.w(w20_78),.acc(r20_78),.res(r20_79),.clk(clk),.wout(w20_79));
	PE pe20_80(.x(x80),.w(w20_79),.acc(r20_79),.res(r20_80),.clk(clk),.wout(w20_80));
	PE pe20_81(.x(x81),.w(w20_80),.acc(r20_80),.res(r20_81),.clk(clk),.wout(w20_81));
	PE pe20_82(.x(x82),.w(w20_81),.acc(r20_81),.res(r20_82),.clk(clk),.wout(w20_82));
	PE pe20_83(.x(x83),.w(w20_82),.acc(r20_82),.res(r20_83),.clk(clk),.wout(w20_83));
	PE pe20_84(.x(x84),.w(w20_83),.acc(r20_83),.res(r20_84),.clk(clk),.wout(w20_84));
	PE pe20_85(.x(x85),.w(w20_84),.acc(r20_84),.res(r20_85),.clk(clk),.wout(w20_85));
	PE pe20_86(.x(x86),.w(w20_85),.acc(r20_85),.res(r20_86),.clk(clk),.wout(w20_86));
	PE pe20_87(.x(x87),.w(w20_86),.acc(r20_86),.res(r20_87),.clk(clk),.wout(w20_87));
	PE pe20_88(.x(x88),.w(w20_87),.acc(r20_87),.res(r20_88),.clk(clk),.wout(w20_88));
	PE pe20_89(.x(x89),.w(w20_88),.acc(r20_88),.res(r20_89),.clk(clk),.wout(w20_89));
	PE pe20_90(.x(x90),.w(w20_89),.acc(r20_89),.res(r20_90),.clk(clk),.wout(w20_90));
	PE pe20_91(.x(x91),.w(w20_90),.acc(r20_90),.res(r20_91),.clk(clk),.wout(w20_91));
	PE pe20_92(.x(x92),.w(w20_91),.acc(r20_91),.res(r20_92),.clk(clk),.wout(w20_92));
	PE pe20_93(.x(x93),.w(w20_92),.acc(r20_92),.res(r20_93),.clk(clk),.wout(w20_93));
	PE pe20_94(.x(x94),.w(w20_93),.acc(r20_93),.res(r20_94),.clk(clk),.wout(w20_94));
	PE pe20_95(.x(x95),.w(w20_94),.acc(r20_94),.res(r20_95),.clk(clk),.wout(w20_95));
	PE pe20_96(.x(x96),.w(w20_95),.acc(r20_95),.res(r20_96),.clk(clk),.wout(w20_96));
	PE pe20_97(.x(x97),.w(w20_96),.acc(r20_96),.res(r20_97),.clk(clk),.wout(w20_97));
	PE pe20_98(.x(x98),.w(w20_97),.acc(r20_97),.res(r20_98),.clk(clk),.wout(w20_98));
	PE pe20_99(.x(x99),.w(w20_98),.acc(r20_98),.res(r20_99),.clk(clk),.wout(w20_99));
	PE pe20_100(.x(x100),.w(w20_99),.acc(r20_99),.res(r20_100),.clk(clk),.wout(w20_100));
	PE pe20_101(.x(x101),.w(w20_100),.acc(r20_100),.res(r20_101),.clk(clk),.wout(w20_101));
	PE pe20_102(.x(x102),.w(w20_101),.acc(r20_101),.res(r20_102),.clk(clk),.wout(w20_102));
	PE pe20_103(.x(x103),.w(w20_102),.acc(r20_102),.res(r20_103),.clk(clk),.wout(w20_103));
	PE pe20_104(.x(x104),.w(w20_103),.acc(r20_103),.res(r20_104),.clk(clk),.wout(w20_104));
	PE pe20_105(.x(x105),.w(w20_104),.acc(r20_104),.res(r20_105),.clk(clk),.wout(w20_105));
	PE pe20_106(.x(x106),.w(w20_105),.acc(r20_105),.res(r20_106),.clk(clk),.wout(w20_106));
	PE pe20_107(.x(x107),.w(w20_106),.acc(r20_106),.res(r20_107),.clk(clk),.wout(w20_107));
	PE pe20_108(.x(x108),.w(w20_107),.acc(r20_107),.res(r20_108),.clk(clk),.wout(w20_108));
	PE pe20_109(.x(x109),.w(w20_108),.acc(r20_108),.res(r20_109),.clk(clk),.wout(w20_109));
	PE pe20_110(.x(x110),.w(w20_109),.acc(r20_109),.res(r20_110),.clk(clk),.wout(w20_110));
	PE pe20_111(.x(x111),.w(w20_110),.acc(r20_110),.res(r20_111),.clk(clk),.wout(w20_111));
	PE pe20_112(.x(x112),.w(w20_111),.acc(r20_111),.res(r20_112),.clk(clk),.wout(w20_112));
	PE pe20_113(.x(x113),.w(w20_112),.acc(r20_112),.res(r20_113),.clk(clk),.wout(w20_113));
	PE pe20_114(.x(x114),.w(w20_113),.acc(r20_113),.res(r20_114),.clk(clk),.wout(w20_114));
	PE pe20_115(.x(x115),.w(w20_114),.acc(r20_114),.res(r20_115),.clk(clk),.wout(w20_115));
	PE pe20_116(.x(x116),.w(w20_115),.acc(r20_115),.res(r20_116),.clk(clk),.wout(w20_116));
	PE pe20_117(.x(x117),.w(w20_116),.acc(r20_116),.res(r20_117),.clk(clk),.wout(w20_117));
	PE pe20_118(.x(x118),.w(w20_117),.acc(r20_117),.res(r20_118),.clk(clk),.wout(w20_118));
	PE pe20_119(.x(x119),.w(w20_118),.acc(r20_118),.res(r20_119),.clk(clk),.wout(w20_119));
	PE pe20_120(.x(x120),.w(w20_119),.acc(r20_119),.res(r20_120),.clk(clk),.wout(w20_120));
	PE pe20_121(.x(x121),.w(w20_120),.acc(r20_120),.res(r20_121),.clk(clk),.wout(w20_121));
	PE pe20_122(.x(x122),.w(w20_121),.acc(r20_121),.res(r20_122),.clk(clk),.wout(w20_122));
	PE pe20_123(.x(x123),.w(w20_122),.acc(r20_122),.res(r20_123),.clk(clk),.wout(w20_123));
	PE pe20_124(.x(x124),.w(w20_123),.acc(r20_123),.res(r20_124),.clk(clk),.wout(w20_124));
	PE pe20_125(.x(x125),.w(w20_124),.acc(r20_124),.res(r20_125),.clk(clk),.wout(w20_125));
	PE pe20_126(.x(x126),.w(w20_125),.acc(r20_125),.res(r20_126),.clk(clk),.wout(w20_126));
	PE pe20_127(.x(x127),.w(w20_126),.acc(r20_126),.res(result20),.clk(clk),.wout(weight20));

	PE pe21_0(.x(x0),.w(w21),.acc(32'h0),.res(r21_0),.clk(clk),.wout(w21_0));
	PE pe21_1(.x(x1),.w(w21_0),.acc(r21_0),.res(r21_1),.clk(clk),.wout(w21_1));
	PE pe21_2(.x(x2),.w(w21_1),.acc(r21_1),.res(r21_2),.clk(clk),.wout(w21_2));
	PE pe21_3(.x(x3),.w(w21_2),.acc(r21_2),.res(r21_3),.clk(clk),.wout(w21_3));
	PE pe21_4(.x(x4),.w(w21_3),.acc(r21_3),.res(r21_4),.clk(clk),.wout(w21_4));
	PE pe21_5(.x(x5),.w(w21_4),.acc(r21_4),.res(r21_5),.clk(clk),.wout(w21_5));
	PE pe21_6(.x(x6),.w(w21_5),.acc(r21_5),.res(r21_6),.clk(clk),.wout(w21_6));
	PE pe21_7(.x(x7),.w(w21_6),.acc(r21_6),.res(r21_7),.clk(clk),.wout(w21_7));
	PE pe21_8(.x(x8),.w(w21_7),.acc(r21_7),.res(r21_8),.clk(clk),.wout(w21_8));
	PE pe21_9(.x(x9),.w(w21_8),.acc(r21_8),.res(r21_9),.clk(clk),.wout(w21_9));
	PE pe21_10(.x(x10),.w(w21_9),.acc(r21_9),.res(r21_10),.clk(clk),.wout(w21_10));
	PE pe21_11(.x(x11),.w(w21_10),.acc(r21_10),.res(r21_11),.clk(clk),.wout(w21_11));
	PE pe21_12(.x(x12),.w(w21_11),.acc(r21_11),.res(r21_12),.clk(clk),.wout(w21_12));
	PE pe21_13(.x(x13),.w(w21_12),.acc(r21_12),.res(r21_13),.clk(clk),.wout(w21_13));
	PE pe21_14(.x(x14),.w(w21_13),.acc(r21_13),.res(r21_14),.clk(clk),.wout(w21_14));
	PE pe21_15(.x(x15),.w(w21_14),.acc(r21_14),.res(r21_15),.clk(clk),.wout(w21_15));
	PE pe21_16(.x(x16),.w(w21_15),.acc(r21_15),.res(r21_16),.clk(clk),.wout(w21_16));
	PE pe21_17(.x(x17),.w(w21_16),.acc(r21_16),.res(r21_17),.clk(clk),.wout(w21_17));
	PE pe21_18(.x(x18),.w(w21_17),.acc(r21_17),.res(r21_18),.clk(clk),.wout(w21_18));
	PE pe21_19(.x(x19),.w(w21_18),.acc(r21_18),.res(r21_19),.clk(clk),.wout(w21_19));
	PE pe21_20(.x(x20),.w(w21_19),.acc(r21_19),.res(r21_20),.clk(clk),.wout(w21_20));
	PE pe21_21(.x(x21),.w(w21_20),.acc(r21_20),.res(r21_21),.clk(clk),.wout(w21_21));
	PE pe21_22(.x(x22),.w(w21_21),.acc(r21_21),.res(r21_22),.clk(clk),.wout(w21_22));
	PE pe21_23(.x(x23),.w(w21_22),.acc(r21_22),.res(r21_23),.clk(clk),.wout(w21_23));
	PE pe21_24(.x(x24),.w(w21_23),.acc(r21_23),.res(r21_24),.clk(clk),.wout(w21_24));
	PE pe21_25(.x(x25),.w(w21_24),.acc(r21_24),.res(r21_25),.clk(clk),.wout(w21_25));
	PE pe21_26(.x(x26),.w(w21_25),.acc(r21_25),.res(r21_26),.clk(clk),.wout(w21_26));
	PE pe21_27(.x(x27),.w(w21_26),.acc(r21_26),.res(r21_27),.clk(clk),.wout(w21_27));
	PE pe21_28(.x(x28),.w(w21_27),.acc(r21_27),.res(r21_28),.clk(clk),.wout(w21_28));
	PE pe21_29(.x(x29),.w(w21_28),.acc(r21_28),.res(r21_29),.clk(clk),.wout(w21_29));
	PE pe21_30(.x(x30),.w(w21_29),.acc(r21_29),.res(r21_30),.clk(clk),.wout(w21_30));
	PE pe21_31(.x(x31),.w(w21_30),.acc(r21_30),.res(r21_31),.clk(clk),.wout(w21_31));
	PE pe21_32(.x(x32),.w(w21_31),.acc(r21_31),.res(r21_32),.clk(clk),.wout(w21_32));
	PE pe21_33(.x(x33),.w(w21_32),.acc(r21_32),.res(r21_33),.clk(clk),.wout(w21_33));
	PE pe21_34(.x(x34),.w(w21_33),.acc(r21_33),.res(r21_34),.clk(clk),.wout(w21_34));
	PE pe21_35(.x(x35),.w(w21_34),.acc(r21_34),.res(r21_35),.clk(clk),.wout(w21_35));
	PE pe21_36(.x(x36),.w(w21_35),.acc(r21_35),.res(r21_36),.clk(clk),.wout(w21_36));
	PE pe21_37(.x(x37),.w(w21_36),.acc(r21_36),.res(r21_37),.clk(clk),.wout(w21_37));
	PE pe21_38(.x(x38),.w(w21_37),.acc(r21_37),.res(r21_38),.clk(clk),.wout(w21_38));
	PE pe21_39(.x(x39),.w(w21_38),.acc(r21_38),.res(r21_39),.clk(clk),.wout(w21_39));
	PE pe21_40(.x(x40),.w(w21_39),.acc(r21_39),.res(r21_40),.clk(clk),.wout(w21_40));
	PE pe21_41(.x(x41),.w(w21_40),.acc(r21_40),.res(r21_41),.clk(clk),.wout(w21_41));
	PE pe21_42(.x(x42),.w(w21_41),.acc(r21_41),.res(r21_42),.clk(clk),.wout(w21_42));
	PE pe21_43(.x(x43),.w(w21_42),.acc(r21_42),.res(r21_43),.clk(clk),.wout(w21_43));
	PE pe21_44(.x(x44),.w(w21_43),.acc(r21_43),.res(r21_44),.clk(clk),.wout(w21_44));
	PE pe21_45(.x(x45),.w(w21_44),.acc(r21_44),.res(r21_45),.clk(clk),.wout(w21_45));
	PE pe21_46(.x(x46),.w(w21_45),.acc(r21_45),.res(r21_46),.clk(clk),.wout(w21_46));
	PE pe21_47(.x(x47),.w(w21_46),.acc(r21_46),.res(r21_47),.clk(clk),.wout(w21_47));
	PE pe21_48(.x(x48),.w(w21_47),.acc(r21_47),.res(r21_48),.clk(clk),.wout(w21_48));
	PE pe21_49(.x(x49),.w(w21_48),.acc(r21_48),.res(r21_49),.clk(clk),.wout(w21_49));
	PE pe21_50(.x(x50),.w(w21_49),.acc(r21_49),.res(r21_50),.clk(clk),.wout(w21_50));
	PE pe21_51(.x(x51),.w(w21_50),.acc(r21_50),.res(r21_51),.clk(clk),.wout(w21_51));
	PE pe21_52(.x(x52),.w(w21_51),.acc(r21_51),.res(r21_52),.clk(clk),.wout(w21_52));
	PE pe21_53(.x(x53),.w(w21_52),.acc(r21_52),.res(r21_53),.clk(clk),.wout(w21_53));
	PE pe21_54(.x(x54),.w(w21_53),.acc(r21_53),.res(r21_54),.clk(clk),.wout(w21_54));
	PE pe21_55(.x(x55),.w(w21_54),.acc(r21_54),.res(r21_55),.clk(clk),.wout(w21_55));
	PE pe21_56(.x(x56),.w(w21_55),.acc(r21_55),.res(r21_56),.clk(clk),.wout(w21_56));
	PE pe21_57(.x(x57),.w(w21_56),.acc(r21_56),.res(r21_57),.clk(clk),.wout(w21_57));
	PE pe21_58(.x(x58),.w(w21_57),.acc(r21_57),.res(r21_58),.clk(clk),.wout(w21_58));
	PE pe21_59(.x(x59),.w(w21_58),.acc(r21_58),.res(r21_59),.clk(clk),.wout(w21_59));
	PE pe21_60(.x(x60),.w(w21_59),.acc(r21_59),.res(r21_60),.clk(clk),.wout(w21_60));
	PE pe21_61(.x(x61),.w(w21_60),.acc(r21_60),.res(r21_61),.clk(clk),.wout(w21_61));
	PE pe21_62(.x(x62),.w(w21_61),.acc(r21_61),.res(r21_62),.clk(clk),.wout(w21_62));
	PE pe21_63(.x(x63),.w(w21_62),.acc(r21_62),.res(r21_63),.clk(clk),.wout(w21_63));
	PE pe21_64(.x(x64),.w(w21_63),.acc(r21_63),.res(r21_64),.clk(clk),.wout(w21_64));
	PE pe21_65(.x(x65),.w(w21_64),.acc(r21_64),.res(r21_65),.clk(clk),.wout(w21_65));
	PE pe21_66(.x(x66),.w(w21_65),.acc(r21_65),.res(r21_66),.clk(clk),.wout(w21_66));
	PE pe21_67(.x(x67),.w(w21_66),.acc(r21_66),.res(r21_67),.clk(clk),.wout(w21_67));
	PE pe21_68(.x(x68),.w(w21_67),.acc(r21_67),.res(r21_68),.clk(clk),.wout(w21_68));
	PE pe21_69(.x(x69),.w(w21_68),.acc(r21_68),.res(r21_69),.clk(clk),.wout(w21_69));
	PE pe21_70(.x(x70),.w(w21_69),.acc(r21_69),.res(r21_70),.clk(clk),.wout(w21_70));
	PE pe21_71(.x(x71),.w(w21_70),.acc(r21_70),.res(r21_71),.clk(clk),.wout(w21_71));
	PE pe21_72(.x(x72),.w(w21_71),.acc(r21_71),.res(r21_72),.clk(clk),.wout(w21_72));
	PE pe21_73(.x(x73),.w(w21_72),.acc(r21_72),.res(r21_73),.clk(clk),.wout(w21_73));
	PE pe21_74(.x(x74),.w(w21_73),.acc(r21_73),.res(r21_74),.clk(clk),.wout(w21_74));
	PE pe21_75(.x(x75),.w(w21_74),.acc(r21_74),.res(r21_75),.clk(clk),.wout(w21_75));
	PE pe21_76(.x(x76),.w(w21_75),.acc(r21_75),.res(r21_76),.clk(clk),.wout(w21_76));
	PE pe21_77(.x(x77),.w(w21_76),.acc(r21_76),.res(r21_77),.clk(clk),.wout(w21_77));
	PE pe21_78(.x(x78),.w(w21_77),.acc(r21_77),.res(r21_78),.clk(clk),.wout(w21_78));
	PE pe21_79(.x(x79),.w(w21_78),.acc(r21_78),.res(r21_79),.clk(clk),.wout(w21_79));
	PE pe21_80(.x(x80),.w(w21_79),.acc(r21_79),.res(r21_80),.clk(clk),.wout(w21_80));
	PE pe21_81(.x(x81),.w(w21_80),.acc(r21_80),.res(r21_81),.clk(clk),.wout(w21_81));
	PE pe21_82(.x(x82),.w(w21_81),.acc(r21_81),.res(r21_82),.clk(clk),.wout(w21_82));
	PE pe21_83(.x(x83),.w(w21_82),.acc(r21_82),.res(r21_83),.clk(clk),.wout(w21_83));
	PE pe21_84(.x(x84),.w(w21_83),.acc(r21_83),.res(r21_84),.clk(clk),.wout(w21_84));
	PE pe21_85(.x(x85),.w(w21_84),.acc(r21_84),.res(r21_85),.clk(clk),.wout(w21_85));
	PE pe21_86(.x(x86),.w(w21_85),.acc(r21_85),.res(r21_86),.clk(clk),.wout(w21_86));
	PE pe21_87(.x(x87),.w(w21_86),.acc(r21_86),.res(r21_87),.clk(clk),.wout(w21_87));
	PE pe21_88(.x(x88),.w(w21_87),.acc(r21_87),.res(r21_88),.clk(clk),.wout(w21_88));
	PE pe21_89(.x(x89),.w(w21_88),.acc(r21_88),.res(r21_89),.clk(clk),.wout(w21_89));
	PE pe21_90(.x(x90),.w(w21_89),.acc(r21_89),.res(r21_90),.clk(clk),.wout(w21_90));
	PE pe21_91(.x(x91),.w(w21_90),.acc(r21_90),.res(r21_91),.clk(clk),.wout(w21_91));
	PE pe21_92(.x(x92),.w(w21_91),.acc(r21_91),.res(r21_92),.clk(clk),.wout(w21_92));
	PE pe21_93(.x(x93),.w(w21_92),.acc(r21_92),.res(r21_93),.clk(clk),.wout(w21_93));
	PE pe21_94(.x(x94),.w(w21_93),.acc(r21_93),.res(r21_94),.clk(clk),.wout(w21_94));
	PE pe21_95(.x(x95),.w(w21_94),.acc(r21_94),.res(r21_95),.clk(clk),.wout(w21_95));
	PE pe21_96(.x(x96),.w(w21_95),.acc(r21_95),.res(r21_96),.clk(clk),.wout(w21_96));
	PE pe21_97(.x(x97),.w(w21_96),.acc(r21_96),.res(r21_97),.clk(clk),.wout(w21_97));
	PE pe21_98(.x(x98),.w(w21_97),.acc(r21_97),.res(r21_98),.clk(clk),.wout(w21_98));
	PE pe21_99(.x(x99),.w(w21_98),.acc(r21_98),.res(r21_99),.clk(clk),.wout(w21_99));
	PE pe21_100(.x(x100),.w(w21_99),.acc(r21_99),.res(r21_100),.clk(clk),.wout(w21_100));
	PE pe21_101(.x(x101),.w(w21_100),.acc(r21_100),.res(r21_101),.clk(clk),.wout(w21_101));
	PE pe21_102(.x(x102),.w(w21_101),.acc(r21_101),.res(r21_102),.clk(clk),.wout(w21_102));
	PE pe21_103(.x(x103),.w(w21_102),.acc(r21_102),.res(r21_103),.clk(clk),.wout(w21_103));
	PE pe21_104(.x(x104),.w(w21_103),.acc(r21_103),.res(r21_104),.clk(clk),.wout(w21_104));
	PE pe21_105(.x(x105),.w(w21_104),.acc(r21_104),.res(r21_105),.clk(clk),.wout(w21_105));
	PE pe21_106(.x(x106),.w(w21_105),.acc(r21_105),.res(r21_106),.clk(clk),.wout(w21_106));
	PE pe21_107(.x(x107),.w(w21_106),.acc(r21_106),.res(r21_107),.clk(clk),.wout(w21_107));
	PE pe21_108(.x(x108),.w(w21_107),.acc(r21_107),.res(r21_108),.clk(clk),.wout(w21_108));
	PE pe21_109(.x(x109),.w(w21_108),.acc(r21_108),.res(r21_109),.clk(clk),.wout(w21_109));
	PE pe21_110(.x(x110),.w(w21_109),.acc(r21_109),.res(r21_110),.clk(clk),.wout(w21_110));
	PE pe21_111(.x(x111),.w(w21_110),.acc(r21_110),.res(r21_111),.clk(clk),.wout(w21_111));
	PE pe21_112(.x(x112),.w(w21_111),.acc(r21_111),.res(r21_112),.clk(clk),.wout(w21_112));
	PE pe21_113(.x(x113),.w(w21_112),.acc(r21_112),.res(r21_113),.clk(clk),.wout(w21_113));
	PE pe21_114(.x(x114),.w(w21_113),.acc(r21_113),.res(r21_114),.clk(clk),.wout(w21_114));
	PE pe21_115(.x(x115),.w(w21_114),.acc(r21_114),.res(r21_115),.clk(clk),.wout(w21_115));
	PE pe21_116(.x(x116),.w(w21_115),.acc(r21_115),.res(r21_116),.clk(clk),.wout(w21_116));
	PE pe21_117(.x(x117),.w(w21_116),.acc(r21_116),.res(r21_117),.clk(clk),.wout(w21_117));
	PE pe21_118(.x(x118),.w(w21_117),.acc(r21_117),.res(r21_118),.clk(clk),.wout(w21_118));
	PE pe21_119(.x(x119),.w(w21_118),.acc(r21_118),.res(r21_119),.clk(clk),.wout(w21_119));
	PE pe21_120(.x(x120),.w(w21_119),.acc(r21_119),.res(r21_120),.clk(clk),.wout(w21_120));
	PE pe21_121(.x(x121),.w(w21_120),.acc(r21_120),.res(r21_121),.clk(clk),.wout(w21_121));
	PE pe21_122(.x(x122),.w(w21_121),.acc(r21_121),.res(r21_122),.clk(clk),.wout(w21_122));
	PE pe21_123(.x(x123),.w(w21_122),.acc(r21_122),.res(r21_123),.clk(clk),.wout(w21_123));
	PE pe21_124(.x(x124),.w(w21_123),.acc(r21_123),.res(r21_124),.clk(clk),.wout(w21_124));
	PE pe21_125(.x(x125),.w(w21_124),.acc(r21_124),.res(r21_125),.clk(clk),.wout(w21_125));
	PE pe21_126(.x(x126),.w(w21_125),.acc(r21_125),.res(r21_126),.clk(clk),.wout(w21_126));
	PE pe21_127(.x(x127),.w(w21_126),.acc(r21_126),.res(result21),.clk(clk),.wout(weight21));

	PE pe22_0(.x(x0),.w(w22),.acc(32'h0),.res(r22_0),.clk(clk),.wout(w22_0));
	PE pe22_1(.x(x1),.w(w22_0),.acc(r22_0),.res(r22_1),.clk(clk),.wout(w22_1));
	PE pe22_2(.x(x2),.w(w22_1),.acc(r22_1),.res(r22_2),.clk(clk),.wout(w22_2));
	PE pe22_3(.x(x3),.w(w22_2),.acc(r22_2),.res(r22_3),.clk(clk),.wout(w22_3));
	PE pe22_4(.x(x4),.w(w22_3),.acc(r22_3),.res(r22_4),.clk(clk),.wout(w22_4));
	PE pe22_5(.x(x5),.w(w22_4),.acc(r22_4),.res(r22_5),.clk(clk),.wout(w22_5));
	PE pe22_6(.x(x6),.w(w22_5),.acc(r22_5),.res(r22_6),.clk(clk),.wout(w22_6));
	PE pe22_7(.x(x7),.w(w22_6),.acc(r22_6),.res(r22_7),.clk(clk),.wout(w22_7));
	PE pe22_8(.x(x8),.w(w22_7),.acc(r22_7),.res(r22_8),.clk(clk),.wout(w22_8));
	PE pe22_9(.x(x9),.w(w22_8),.acc(r22_8),.res(r22_9),.clk(clk),.wout(w22_9));
	PE pe22_10(.x(x10),.w(w22_9),.acc(r22_9),.res(r22_10),.clk(clk),.wout(w22_10));
	PE pe22_11(.x(x11),.w(w22_10),.acc(r22_10),.res(r22_11),.clk(clk),.wout(w22_11));
	PE pe22_12(.x(x12),.w(w22_11),.acc(r22_11),.res(r22_12),.clk(clk),.wout(w22_12));
	PE pe22_13(.x(x13),.w(w22_12),.acc(r22_12),.res(r22_13),.clk(clk),.wout(w22_13));
	PE pe22_14(.x(x14),.w(w22_13),.acc(r22_13),.res(r22_14),.clk(clk),.wout(w22_14));
	PE pe22_15(.x(x15),.w(w22_14),.acc(r22_14),.res(r22_15),.clk(clk),.wout(w22_15));
	PE pe22_16(.x(x16),.w(w22_15),.acc(r22_15),.res(r22_16),.clk(clk),.wout(w22_16));
	PE pe22_17(.x(x17),.w(w22_16),.acc(r22_16),.res(r22_17),.clk(clk),.wout(w22_17));
	PE pe22_18(.x(x18),.w(w22_17),.acc(r22_17),.res(r22_18),.clk(clk),.wout(w22_18));
	PE pe22_19(.x(x19),.w(w22_18),.acc(r22_18),.res(r22_19),.clk(clk),.wout(w22_19));
	PE pe22_20(.x(x20),.w(w22_19),.acc(r22_19),.res(r22_20),.clk(clk),.wout(w22_20));
	PE pe22_21(.x(x21),.w(w22_20),.acc(r22_20),.res(r22_21),.clk(clk),.wout(w22_21));
	PE pe22_22(.x(x22),.w(w22_21),.acc(r22_21),.res(r22_22),.clk(clk),.wout(w22_22));
	PE pe22_23(.x(x23),.w(w22_22),.acc(r22_22),.res(r22_23),.clk(clk),.wout(w22_23));
	PE pe22_24(.x(x24),.w(w22_23),.acc(r22_23),.res(r22_24),.clk(clk),.wout(w22_24));
	PE pe22_25(.x(x25),.w(w22_24),.acc(r22_24),.res(r22_25),.clk(clk),.wout(w22_25));
	PE pe22_26(.x(x26),.w(w22_25),.acc(r22_25),.res(r22_26),.clk(clk),.wout(w22_26));
	PE pe22_27(.x(x27),.w(w22_26),.acc(r22_26),.res(r22_27),.clk(clk),.wout(w22_27));
	PE pe22_28(.x(x28),.w(w22_27),.acc(r22_27),.res(r22_28),.clk(clk),.wout(w22_28));
	PE pe22_29(.x(x29),.w(w22_28),.acc(r22_28),.res(r22_29),.clk(clk),.wout(w22_29));
	PE pe22_30(.x(x30),.w(w22_29),.acc(r22_29),.res(r22_30),.clk(clk),.wout(w22_30));
	PE pe22_31(.x(x31),.w(w22_30),.acc(r22_30),.res(r22_31),.clk(clk),.wout(w22_31));
	PE pe22_32(.x(x32),.w(w22_31),.acc(r22_31),.res(r22_32),.clk(clk),.wout(w22_32));
	PE pe22_33(.x(x33),.w(w22_32),.acc(r22_32),.res(r22_33),.clk(clk),.wout(w22_33));
	PE pe22_34(.x(x34),.w(w22_33),.acc(r22_33),.res(r22_34),.clk(clk),.wout(w22_34));
	PE pe22_35(.x(x35),.w(w22_34),.acc(r22_34),.res(r22_35),.clk(clk),.wout(w22_35));
	PE pe22_36(.x(x36),.w(w22_35),.acc(r22_35),.res(r22_36),.clk(clk),.wout(w22_36));
	PE pe22_37(.x(x37),.w(w22_36),.acc(r22_36),.res(r22_37),.clk(clk),.wout(w22_37));
	PE pe22_38(.x(x38),.w(w22_37),.acc(r22_37),.res(r22_38),.clk(clk),.wout(w22_38));
	PE pe22_39(.x(x39),.w(w22_38),.acc(r22_38),.res(r22_39),.clk(clk),.wout(w22_39));
	PE pe22_40(.x(x40),.w(w22_39),.acc(r22_39),.res(r22_40),.clk(clk),.wout(w22_40));
	PE pe22_41(.x(x41),.w(w22_40),.acc(r22_40),.res(r22_41),.clk(clk),.wout(w22_41));
	PE pe22_42(.x(x42),.w(w22_41),.acc(r22_41),.res(r22_42),.clk(clk),.wout(w22_42));
	PE pe22_43(.x(x43),.w(w22_42),.acc(r22_42),.res(r22_43),.clk(clk),.wout(w22_43));
	PE pe22_44(.x(x44),.w(w22_43),.acc(r22_43),.res(r22_44),.clk(clk),.wout(w22_44));
	PE pe22_45(.x(x45),.w(w22_44),.acc(r22_44),.res(r22_45),.clk(clk),.wout(w22_45));
	PE pe22_46(.x(x46),.w(w22_45),.acc(r22_45),.res(r22_46),.clk(clk),.wout(w22_46));
	PE pe22_47(.x(x47),.w(w22_46),.acc(r22_46),.res(r22_47),.clk(clk),.wout(w22_47));
	PE pe22_48(.x(x48),.w(w22_47),.acc(r22_47),.res(r22_48),.clk(clk),.wout(w22_48));
	PE pe22_49(.x(x49),.w(w22_48),.acc(r22_48),.res(r22_49),.clk(clk),.wout(w22_49));
	PE pe22_50(.x(x50),.w(w22_49),.acc(r22_49),.res(r22_50),.clk(clk),.wout(w22_50));
	PE pe22_51(.x(x51),.w(w22_50),.acc(r22_50),.res(r22_51),.clk(clk),.wout(w22_51));
	PE pe22_52(.x(x52),.w(w22_51),.acc(r22_51),.res(r22_52),.clk(clk),.wout(w22_52));
	PE pe22_53(.x(x53),.w(w22_52),.acc(r22_52),.res(r22_53),.clk(clk),.wout(w22_53));
	PE pe22_54(.x(x54),.w(w22_53),.acc(r22_53),.res(r22_54),.clk(clk),.wout(w22_54));
	PE pe22_55(.x(x55),.w(w22_54),.acc(r22_54),.res(r22_55),.clk(clk),.wout(w22_55));
	PE pe22_56(.x(x56),.w(w22_55),.acc(r22_55),.res(r22_56),.clk(clk),.wout(w22_56));
	PE pe22_57(.x(x57),.w(w22_56),.acc(r22_56),.res(r22_57),.clk(clk),.wout(w22_57));
	PE pe22_58(.x(x58),.w(w22_57),.acc(r22_57),.res(r22_58),.clk(clk),.wout(w22_58));
	PE pe22_59(.x(x59),.w(w22_58),.acc(r22_58),.res(r22_59),.clk(clk),.wout(w22_59));
	PE pe22_60(.x(x60),.w(w22_59),.acc(r22_59),.res(r22_60),.clk(clk),.wout(w22_60));
	PE pe22_61(.x(x61),.w(w22_60),.acc(r22_60),.res(r22_61),.clk(clk),.wout(w22_61));
	PE pe22_62(.x(x62),.w(w22_61),.acc(r22_61),.res(r22_62),.clk(clk),.wout(w22_62));
	PE pe22_63(.x(x63),.w(w22_62),.acc(r22_62),.res(r22_63),.clk(clk),.wout(w22_63));
	PE pe22_64(.x(x64),.w(w22_63),.acc(r22_63),.res(r22_64),.clk(clk),.wout(w22_64));
	PE pe22_65(.x(x65),.w(w22_64),.acc(r22_64),.res(r22_65),.clk(clk),.wout(w22_65));
	PE pe22_66(.x(x66),.w(w22_65),.acc(r22_65),.res(r22_66),.clk(clk),.wout(w22_66));
	PE pe22_67(.x(x67),.w(w22_66),.acc(r22_66),.res(r22_67),.clk(clk),.wout(w22_67));
	PE pe22_68(.x(x68),.w(w22_67),.acc(r22_67),.res(r22_68),.clk(clk),.wout(w22_68));
	PE pe22_69(.x(x69),.w(w22_68),.acc(r22_68),.res(r22_69),.clk(clk),.wout(w22_69));
	PE pe22_70(.x(x70),.w(w22_69),.acc(r22_69),.res(r22_70),.clk(clk),.wout(w22_70));
	PE pe22_71(.x(x71),.w(w22_70),.acc(r22_70),.res(r22_71),.clk(clk),.wout(w22_71));
	PE pe22_72(.x(x72),.w(w22_71),.acc(r22_71),.res(r22_72),.clk(clk),.wout(w22_72));
	PE pe22_73(.x(x73),.w(w22_72),.acc(r22_72),.res(r22_73),.clk(clk),.wout(w22_73));
	PE pe22_74(.x(x74),.w(w22_73),.acc(r22_73),.res(r22_74),.clk(clk),.wout(w22_74));
	PE pe22_75(.x(x75),.w(w22_74),.acc(r22_74),.res(r22_75),.clk(clk),.wout(w22_75));
	PE pe22_76(.x(x76),.w(w22_75),.acc(r22_75),.res(r22_76),.clk(clk),.wout(w22_76));
	PE pe22_77(.x(x77),.w(w22_76),.acc(r22_76),.res(r22_77),.clk(clk),.wout(w22_77));
	PE pe22_78(.x(x78),.w(w22_77),.acc(r22_77),.res(r22_78),.clk(clk),.wout(w22_78));
	PE pe22_79(.x(x79),.w(w22_78),.acc(r22_78),.res(r22_79),.clk(clk),.wout(w22_79));
	PE pe22_80(.x(x80),.w(w22_79),.acc(r22_79),.res(r22_80),.clk(clk),.wout(w22_80));
	PE pe22_81(.x(x81),.w(w22_80),.acc(r22_80),.res(r22_81),.clk(clk),.wout(w22_81));
	PE pe22_82(.x(x82),.w(w22_81),.acc(r22_81),.res(r22_82),.clk(clk),.wout(w22_82));
	PE pe22_83(.x(x83),.w(w22_82),.acc(r22_82),.res(r22_83),.clk(clk),.wout(w22_83));
	PE pe22_84(.x(x84),.w(w22_83),.acc(r22_83),.res(r22_84),.clk(clk),.wout(w22_84));
	PE pe22_85(.x(x85),.w(w22_84),.acc(r22_84),.res(r22_85),.clk(clk),.wout(w22_85));
	PE pe22_86(.x(x86),.w(w22_85),.acc(r22_85),.res(r22_86),.clk(clk),.wout(w22_86));
	PE pe22_87(.x(x87),.w(w22_86),.acc(r22_86),.res(r22_87),.clk(clk),.wout(w22_87));
	PE pe22_88(.x(x88),.w(w22_87),.acc(r22_87),.res(r22_88),.clk(clk),.wout(w22_88));
	PE pe22_89(.x(x89),.w(w22_88),.acc(r22_88),.res(r22_89),.clk(clk),.wout(w22_89));
	PE pe22_90(.x(x90),.w(w22_89),.acc(r22_89),.res(r22_90),.clk(clk),.wout(w22_90));
	PE pe22_91(.x(x91),.w(w22_90),.acc(r22_90),.res(r22_91),.clk(clk),.wout(w22_91));
	PE pe22_92(.x(x92),.w(w22_91),.acc(r22_91),.res(r22_92),.clk(clk),.wout(w22_92));
	PE pe22_93(.x(x93),.w(w22_92),.acc(r22_92),.res(r22_93),.clk(clk),.wout(w22_93));
	PE pe22_94(.x(x94),.w(w22_93),.acc(r22_93),.res(r22_94),.clk(clk),.wout(w22_94));
	PE pe22_95(.x(x95),.w(w22_94),.acc(r22_94),.res(r22_95),.clk(clk),.wout(w22_95));
	PE pe22_96(.x(x96),.w(w22_95),.acc(r22_95),.res(r22_96),.clk(clk),.wout(w22_96));
	PE pe22_97(.x(x97),.w(w22_96),.acc(r22_96),.res(r22_97),.clk(clk),.wout(w22_97));
	PE pe22_98(.x(x98),.w(w22_97),.acc(r22_97),.res(r22_98),.clk(clk),.wout(w22_98));
	PE pe22_99(.x(x99),.w(w22_98),.acc(r22_98),.res(r22_99),.clk(clk),.wout(w22_99));
	PE pe22_100(.x(x100),.w(w22_99),.acc(r22_99),.res(r22_100),.clk(clk),.wout(w22_100));
	PE pe22_101(.x(x101),.w(w22_100),.acc(r22_100),.res(r22_101),.clk(clk),.wout(w22_101));
	PE pe22_102(.x(x102),.w(w22_101),.acc(r22_101),.res(r22_102),.clk(clk),.wout(w22_102));
	PE pe22_103(.x(x103),.w(w22_102),.acc(r22_102),.res(r22_103),.clk(clk),.wout(w22_103));
	PE pe22_104(.x(x104),.w(w22_103),.acc(r22_103),.res(r22_104),.clk(clk),.wout(w22_104));
	PE pe22_105(.x(x105),.w(w22_104),.acc(r22_104),.res(r22_105),.clk(clk),.wout(w22_105));
	PE pe22_106(.x(x106),.w(w22_105),.acc(r22_105),.res(r22_106),.clk(clk),.wout(w22_106));
	PE pe22_107(.x(x107),.w(w22_106),.acc(r22_106),.res(r22_107),.clk(clk),.wout(w22_107));
	PE pe22_108(.x(x108),.w(w22_107),.acc(r22_107),.res(r22_108),.clk(clk),.wout(w22_108));
	PE pe22_109(.x(x109),.w(w22_108),.acc(r22_108),.res(r22_109),.clk(clk),.wout(w22_109));
	PE pe22_110(.x(x110),.w(w22_109),.acc(r22_109),.res(r22_110),.clk(clk),.wout(w22_110));
	PE pe22_111(.x(x111),.w(w22_110),.acc(r22_110),.res(r22_111),.clk(clk),.wout(w22_111));
	PE pe22_112(.x(x112),.w(w22_111),.acc(r22_111),.res(r22_112),.clk(clk),.wout(w22_112));
	PE pe22_113(.x(x113),.w(w22_112),.acc(r22_112),.res(r22_113),.clk(clk),.wout(w22_113));
	PE pe22_114(.x(x114),.w(w22_113),.acc(r22_113),.res(r22_114),.clk(clk),.wout(w22_114));
	PE pe22_115(.x(x115),.w(w22_114),.acc(r22_114),.res(r22_115),.clk(clk),.wout(w22_115));
	PE pe22_116(.x(x116),.w(w22_115),.acc(r22_115),.res(r22_116),.clk(clk),.wout(w22_116));
	PE pe22_117(.x(x117),.w(w22_116),.acc(r22_116),.res(r22_117),.clk(clk),.wout(w22_117));
	PE pe22_118(.x(x118),.w(w22_117),.acc(r22_117),.res(r22_118),.clk(clk),.wout(w22_118));
	PE pe22_119(.x(x119),.w(w22_118),.acc(r22_118),.res(r22_119),.clk(clk),.wout(w22_119));
	PE pe22_120(.x(x120),.w(w22_119),.acc(r22_119),.res(r22_120),.clk(clk),.wout(w22_120));
	PE pe22_121(.x(x121),.w(w22_120),.acc(r22_120),.res(r22_121),.clk(clk),.wout(w22_121));
	PE pe22_122(.x(x122),.w(w22_121),.acc(r22_121),.res(r22_122),.clk(clk),.wout(w22_122));
	PE pe22_123(.x(x123),.w(w22_122),.acc(r22_122),.res(r22_123),.clk(clk),.wout(w22_123));
	PE pe22_124(.x(x124),.w(w22_123),.acc(r22_123),.res(r22_124),.clk(clk),.wout(w22_124));
	PE pe22_125(.x(x125),.w(w22_124),.acc(r22_124),.res(r22_125),.clk(clk),.wout(w22_125));
	PE pe22_126(.x(x126),.w(w22_125),.acc(r22_125),.res(r22_126),.clk(clk),.wout(w22_126));
	PE pe22_127(.x(x127),.w(w22_126),.acc(r22_126),.res(result22),.clk(clk),.wout(weight22));

	PE pe23_0(.x(x0),.w(w23),.acc(32'h0),.res(r23_0),.clk(clk),.wout(w23_0));
	PE pe23_1(.x(x1),.w(w23_0),.acc(r23_0),.res(r23_1),.clk(clk),.wout(w23_1));
	PE pe23_2(.x(x2),.w(w23_1),.acc(r23_1),.res(r23_2),.clk(clk),.wout(w23_2));
	PE pe23_3(.x(x3),.w(w23_2),.acc(r23_2),.res(r23_3),.clk(clk),.wout(w23_3));
	PE pe23_4(.x(x4),.w(w23_3),.acc(r23_3),.res(r23_4),.clk(clk),.wout(w23_4));
	PE pe23_5(.x(x5),.w(w23_4),.acc(r23_4),.res(r23_5),.clk(clk),.wout(w23_5));
	PE pe23_6(.x(x6),.w(w23_5),.acc(r23_5),.res(r23_6),.clk(clk),.wout(w23_6));
	PE pe23_7(.x(x7),.w(w23_6),.acc(r23_6),.res(r23_7),.clk(clk),.wout(w23_7));
	PE pe23_8(.x(x8),.w(w23_7),.acc(r23_7),.res(r23_8),.clk(clk),.wout(w23_8));
	PE pe23_9(.x(x9),.w(w23_8),.acc(r23_8),.res(r23_9),.clk(clk),.wout(w23_9));
	PE pe23_10(.x(x10),.w(w23_9),.acc(r23_9),.res(r23_10),.clk(clk),.wout(w23_10));
	PE pe23_11(.x(x11),.w(w23_10),.acc(r23_10),.res(r23_11),.clk(clk),.wout(w23_11));
	PE pe23_12(.x(x12),.w(w23_11),.acc(r23_11),.res(r23_12),.clk(clk),.wout(w23_12));
	PE pe23_13(.x(x13),.w(w23_12),.acc(r23_12),.res(r23_13),.clk(clk),.wout(w23_13));
	PE pe23_14(.x(x14),.w(w23_13),.acc(r23_13),.res(r23_14),.clk(clk),.wout(w23_14));
	PE pe23_15(.x(x15),.w(w23_14),.acc(r23_14),.res(r23_15),.clk(clk),.wout(w23_15));
	PE pe23_16(.x(x16),.w(w23_15),.acc(r23_15),.res(r23_16),.clk(clk),.wout(w23_16));
	PE pe23_17(.x(x17),.w(w23_16),.acc(r23_16),.res(r23_17),.clk(clk),.wout(w23_17));
	PE pe23_18(.x(x18),.w(w23_17),.acc(r23_17),.res(r23_18),.clk(clk),.wout(w23_18));
	PE pe23_19(.x(x19),.w(w23_18),.acc(r23_18),.res(r23_19),.clk(clk),.wout(w23_19));
	PE pe23_20(.x(x20),.w(w23_19),.acc(r23_19),.res(r23_20),.clk(clk),.wout(w23_20));
	PE pe23_21(.x(x21),.w(w23_20),.acc(r23_20),.res(r23_21),.clk(clk),.wout(w23_21));
	PE pe23_22(.x(x22),.w(w23_21),.acc(r23_21),.res(r23_22),.clk(clk),.wout(w23_22));
	PE pe23_23(.x(x23),.w(w23_22),.acc(r23_22),.res(r23_23),.clk(clk),.wout(w23_23));
	PE pe23_24(.x(x24),.w(w23_23),.acc(r23_23),.res(r23_24),.clk(clk),.wout(w23_24));
	PE pe23_25(.x(x25),.w(w23_24),.acc(r23_24),.res(r23_25),.clk(clk),.wout(w23_25));
	PE pe23_26(.x(x26),.w(w23_25),.acc(r23_25),.res(r23_26),.clk(clk),.wout(w23_26));
	PE pe23_27(.x(x27),.w(w23_26),.acc(r23_26),.res(r23_27),.clk(clk),.wout(w23_27));
	PE pe23_28(.x(x28),.w(w23_27),.acc(r23_27),.res(r23_28),.clk(clk),.wout(w23_28));
	PE pe23_29(.x(x29),.w(w23_28),.acc(r23_28),.res(r23_29),.clk(clk),.wout(w23_29));
	PE pe23_30(.x(x30),.w(w23_29),.acc(r23_29),.res(r23_30),.clk(clk),.wout(w23_30));
	PE pe23_31(.x(x31),.w(w23_30),.acc(r23_30),.res(r23_31),.clk(clk),.wout(w23_31));
	PE pe23_32(.x(x32),.w(w23_31),.acc(r23_31),.res(r23_32),.clk(clk),.wout(w23_32));
	PE pe23_33(.x(x33),.w(w23_32),.acc(r23_32),.res(r23_33),.clk(clk),.wout(w23_33));
	PE pe23_34(.x(x34),.w(w23_33),.acc(r23_33),.res(r23_34),.clk(clk),.wout(w23_34));
	PE pe23_35(.x(x35),.w(w23_34),.acc(r23_34),.res(r23_35),.clk(clk),.wout(w23_35));
	PE pe23_36(.x(x36),.w(w23_35),.acc(r23_35),.res(r23_36),.clk(clk),.wout(w23_36));
	PE pe23_37(.x(x37),.w(w23_36),.acc(r23_36),.res(r23_37),.clk(clk),.wout(w23_37));
	PE pe23_38(.x(x38),.w(w23_37),.acc(r23_37),.res(r23_38),.clk(clk),.wout(w23_38));
	PE pe23_39(.x(x39),.w(w23_38),.acc(r23_38),.res(r23_39),.clk(clk),.wout(w23_39));
	PE pe23_40(.x(x40),.w(w23_39),.acc(r23_39),.res(r23_40),.clk(clk),.wout(w23_40));
	PE pe23_41(.x(x41),.w(w23_40),.acc(r23_40),.res(r23_41),.clk(clk),.wout(w23_41));
	PE pe23_42(.x(x42),.w(w23_41),.acc(r23_41),.res(r23_42),.clk(clk),.wout(w23_42));
	PE pe23_43(.x(x43),.w(w23_42),.acc(r23_42),.res(r23_43),.clk(clk),.wout(w23_43));
	PE pe23_44(.x(x44),.w(w23_43),.acc(r23_43),.res(r23_44),.clk(clk),.wout(w23_44));
	PE pe23_45(.x(x45),.w(w23_44),.acc(r23_44),.res(r23_45),.clk(clk),.wout(w23_45));
	PE pe23_46(.x(x46),.w(w23_45),.acc(r23_45),.res(r23_46),.clk(clk),.wout(w23_46));
	PE pe23_47(.x(x47),.w(w23_46),.acc(r23_46),.res(r23_47),.clk(clk),.wout(w23_47));
	PE pe23_48(.x(x48),.w(w23_47),.acc(r23_47),.res(r23_48),.clk(clk),.wout(w23_48));
	PE pe23_49(.x(x49),.w(w23_48),.acc(r23_48),.res(r23_49),.clk(clk),.wout(w23_49));
	PE pe23_50(.x(x50),.w(w23_49),.acc(r23_49),.res(r23_50),.clk(clk),.wout(w23_50));
	PE pe23_51(.x(x51),.w(w23_50),.acc(r23_50),.res(r23_51),.clk(clk),.wout(w23_51));
	PE pe23_52(.x(x52),.w(w23_51),.acc(r23_51),.res(r23_52),.clk(clk),.wout(w23_52));
	PE pe23_53(.x(x53),.w(w23_52),.acc(r23_52),.res(r23_53),.clk(clk),.wout(w23_53));
	PE pe23_54(.x(x54),.w(w23_53),.acc(r23_53),.res(r23_54),.clk(clk),.wout(w23_54));
	PE pe23_55(.x(x55),.w(w23_54),.acc(r23_54),.res(r23_55),.clk(clk),.wout(w23_55));
	PE pe23_56(.x(x56),.w(w23_55),.acc(r23_55),.res(r23_56),.clk(clk),.wout(w23_56));
	PE pe23_57(.x(x57),.w(w23_56),.acc(r23_56),.res(r23_57),.clk(clk),.wout(w23_57));
	PE pe23_58(.x(x58),.w(w23_57),.acc(r23_57),.res(r23_58),.clk(clk),.wout(w23_58));
	PE pe23_59(.x(x59),.w(w23_58),.acc(r23_58),.res(r23_59),.clk(clk),.wout(w23_59));
	PE pe23_60(.x(x60),.w(w23_59),.acc(r23_59),.res(r23_60),.clk(clk),.wout(w23_60));
	PE pe23_61(.x(x61),.w(w23_60),.acc(r23_60),.res(r23_61),.clk(clk),.wout(w23_61));
	PE pe23_62(.x(x62),.w(w23_61),.acc(r23_61),.res(r23_62),.clk(clk),.wout(w23_62));
	PE pe23_63(.x(x63),.w(w23_62),.acc(r23_62),.res(r23_63),.clk(clk),.wout(w23_63));
	PE pe23_64(.x(x64),.w(w23_63),.acc(r23_63),.res(r23_64),.clk(clk),.wout(w23_64));
	PE pe23_65(.x(x65),.w(w23_64),.acc(r23_64),.res(r23_65),.clk(clk),.wout(w23_65));
	PE pe23_66(.x(x66),.w(w23_65),.acc(r23_65),.res(r23_66),.clk(clk),.wout(w23_66));
	PE pe23_67(.x(x67),.w(w23_66),.acc(r23_66),.res(r23_67),.clk(clk),.wout(w23_67));
	PE pe23_68(.x(x68),.w(w23_67),.acc(r23_67),.res(r23_68),.clk(clk),.wout(w23_68));
	PE pe23_69(.x(x69),.w(w23_68),.acc(r23_68),.res(r23_69),.clk(clk),.wout(w23_69));
	PE pe23_70(.x(x70),.w(w23_69),.acc(r23_69),.res(r23_70),.clk(clk),.wout(w23_70));
	PE pe23_71(.x(x71),.w(w23_70),.acc(r23_70),.res(r23_71),.clk(clk),.wout(w23_71));
	PE pe23_72(.x(x72),.w(w23_71),.acc(r23_71),.res(r23_72),.clk(clk),.wout(w23_72));
	PE pe23_73(.x(x73),.w(w23_72),.acc(r23_72),.res(r23_73),.clk(clk),.wout(w23_73));
	PE pe23_74(.x(x74),.w(w23_73),.acc(r23_73),.res(r23_74),.clk(clk),.wout(w23_74));
	PE pe23_75(.x(x75),.w(w23_74),.acc(r23_74),.res(r23_75),.clk(clk),.wout(w23_75));
	PE pe23_76(.x(x76),.w(w23_75),.acc(r23_75),.res(r23_76),.clk(clk),.wout(w23_76));
	PE pe23_77(.x(x77),.w(w23_76),.acc(r23_76),.res(r23_77),.clk(clk),.wout(w23_77));
	PE pe23_78(.x(x78),.w(w23_77),.acc(r23_77),.res(r23_78),.clk(clk),.wout(w23_78));
	PE pe23_79(.x(x79),.w(w23_78),.acc(r23_78),.res(r23_79),.clk(clk),.wout(w23_79));
	PE pe23_80(.x(x80),.w(w23_79),.acc(r23_79),.res(r23_80),.clk(clk),.wout(w23_80));
	PE pe23_81(.x(x81),.w(w23_80),.acc(r23_80),.res(r23_81),.clk(clk),.wout(w23_81));
	PE pe23_82(.x(x82),.w(w23_81),.acc(r23_81),.res(r23_82),.clk(clk),.wout(w23_82));
	PE pe23_83(.x(x83),.w(w23_82),.acc(r23_82),.res(r23_83),.clk(clk),.wout(w23_83));
	PE pe23_84(.x(x84),.w(w23_83),.acc(r23_83),.res(r23_84),.clk(clk),.wout(w23_84));
	PE pe23_85(.x(x85),.w(w23_84),.acc(r23_84),.res(r23_85),.clk(clk),.wout(w23_85));
	PE pe23_86(.x(x86),.w(w23_85),.acc(r23_85),.res(r23_86),.clk(clk),.wout(w23_86));
	PE pe23_87(.x(x87),.w(w23_86),.acc(r23_86),.res(r23_87),.clk(clk),.wout(w23_87));
	PE pe23_88(.x(x88),.w(w23_87),.acc(r23_87),.res(r23_88),.clk(clk),.wout(w23_88));
	PE pe23_89(.x(x89),.w(w23_88),.acc(r23_88),.res(r23_89),.clk(clk),.wout(w23_89));
	PE pe23_90(.x(x90),.w(w23_89),.acc(r23_89),.res(r23_90),.clk(clk),.wout(w23_90));
	PE pe23_91(.x(x91),.w(w23_90),.acc(r23_90),.res(r23_91),.clk(clk),.wout(w23_91));
	PE pe23_92(.x(x92),.w(w23_91),.acc(r23_91),.res(r23_92),.clk(clk),.wout(w23_92));
	PE pe23_93(.x(x93),.w(w23_92),.acc(r23_92),.res(r23_93),.clk(clk),.wout(w23_93));
	PE pe23_94(.x(x94),.w(w23_93),.acc(r23_93),.res(r23_94),.clk(clk),.wout(w23_94));
	PE pe23_95(.x(x95),.w(w23_94),.acc(r23_94),.res(r23_95),.clk(clk),.wout(w23_95));
	PE pe23_96(.x(x96),.w(w23_95),.acc(r23_95),.res(r23_96),.clk(clk),.wout(w23_96));
	PE pe23_97(.x(x97),.w(w23_96),.acc(r23_96),.res(r23_97),.clk(clk),.wout(w23_97));
	PE pe23_98(.x(x98),.w(w23_97),.acc(r23_97),.res(r23_98),.clk(clk),.wout(w23_98));
	PE pe23_99(.x(x99),.w(w23_98),.acc(r23_98),.res(r23_99),.clk(clk),.wout(w23_99));
	PE pe23_100(.x(x100),.w(w23_99),.acc(r23_99),.res(r23_100),.clk(clk),.wout(w23_100));
	PE pe23_101(.x(x101),.w(w23_100),.acc(r23_100),.res(r23_101),.clk(clk),.wout(w23_101));
	PE pe23_102(.x(x102),.w(w23_101),.acc(r23_101),.res(r23_102),.clk(clk),.wout(w23_102));
	PE pe23_103(.x(x103),.w(w23_102),.acc(r23_102),.res(r23_103),.clk(clk),.wout(w23_103));
	PE pe23_104(.x(x104),.w(w23_103),.acc(r23_103),.res(r23_104),.clk(clk),.wout(w23_104));
	PE pe23_105(.x(x105),.w(w23_104),.acc(r23_104),.res(r23_105),.clk(clk),.wout(w23_105));
	PE pe23_106(.x(x106),.w(w23_105),.acc(r23_105),.res(r23_106),.clk(clk),.wout(w23_106));
	PE pe23_107(.x(x107),.w(w23_106),.acc(r23_106),.res(r23_107),.clk(clk),.wout(w23_107));
	PE pe23_108(.x(x108),.w(w23_107),.acc(r23_107),.res(r23_108),.clk(clk),.wout(w23_108));
	PE pe23_109(.x(x109),.w(w23_108),.acc(r23_108),.res(r23_109),.clk(clk),.wout(w23_109));
	PE pe23_110(.x(x110),.w(w23_109),.acc(r23_109),.res(r23_110),.clk(clk),.wout(w23_110));
	PE pe23_111(.x(x111),.w(w23_110),.acc(r23_110),.res(r23_111),.clk(clk),.wout(w23_111));
	PE pe23_112(.x(x112),.w(w23_111),.acc(r23_111),.res(r23_112),.clk(clk),.wout(w23_112));
	PE pe23_113(.x(x113),.w(w23_112),.acc(r23_112),.res(r23_113),.clk(clk),.wout(w23_113));
	PE pe23_114(.x(x114),.w(w23_113),.acc(r23_113),.res(r23_114),.clk(clk),.wout(w23_114));
	PE pe23_115(.x(x115),.w(w23_114),.acc(r23_114),.res(r23_115),.clk(clk),.wout(w23_115));
	PE pe23_116(.x(x116),.w(w23_115),.acc(r23_115),.res(r23_116),.clk(clk),.wout(w23_116));
	PE pe23_117(.x(x117),.w(w23_116),.acc(r23_116),.res(r23_117),.clk(clk),.wout(w23_117));
	PE pe23_118(.x(x118),.w(w23_117),.acc(r23_117),.res(r23_118),.clk(clk),.wout(w23_118));
	PE pe23_119(.x(x119),.w(w23_118),.acc(r23_118),.res(r23_119),.clk(clk),.wout(w23_119));
	PE pe23_120(.x(x120),.w(w23_119),.acc(r23_119),.res(r23_120),.clk(clk),.wout(w23_120));
	PE pe23_121(.x(x121),.w(w23_120),.acc(r23_120),.res(r23_121),.clk(clk),.wout(w23_121));
	PE pe23_122(.x(x122),.w(w23_121),.acc(r23_121),.res(r23_122),.clk(clk),.wout(w23_122));
	PE pe23_123(.x(x123),.w(w23_122),.acc(r23_122),.res(r23_123),.clk(clk),.wout(w23_123));
	PE pe23_124(.x(x124),.w(w23_123),.acc(r23_123),.res(r23_124),.clk(clk),.wout(w23_124));
	PE pe23_125(.x(x125),.w(w23_124),.acc(r23_124),.res(r23_125),.clk(clk),.wout(w23_125));
	PE pe23_126(.x(x126),.w(w23_125),.acc(r23_125),.res(r23_126),.clk(clk),.wout(w23_126));
	PE pe23_127(.x(x127),.w(w23_126),.acc(r23_126),.res(result23),.clk(clk),.wout(weight23));

	PE pe24_0(.x(x0),.w(w24),.acc(32'h0),.res(r24_0),.clk(clk),.wout(w24_0));
	PE pe24_1(.x(x1),.w(w24_0),.acc(r24_0),.res(r24_1),.clk(clk),.wout(w24_1));
	PE pe24_2(.x(x2),.w(w24_1),.acc(r24_1),.res(r24_2),.clk(clk),.wout(w24_2));
	PE pe24_3(.x(x3),.w(w24_2),.acc(r24_2),.res(r24_3),.clk(clk),.wout(w24_3));
	PE pe24_4(.x(x4),.w(w24_3),.acc(r24_3),.res(r24_4),.clk(clk),.wout(w24_4));
	PE pe24_5(.x(x5),.w(w24_4),.acc(r24_4),.res(r24_5),.clk(clk),.wout(w24_5));
	PE pe24_6(.x(x6),.w(w24_5),.acc(r24_5),.res(r24_6),.clk(clk),.wout(w24_6));
	PE pe24_7(.x(x7),.w(w24_6),.acc(r24_6),.res(r24_7),.clk(clk),.wout(w24_7));
	PE pe24_8(.x(x8),.w(w24_7),.acc(r24_7),.res(r24_8),.clk(clk),.wout(w24_8));
	PE pe24_9(.x(x9),.w(w24_8),.acc(r24_8),.res(r24_9),.clk(clk),.wout(w24_9));
	PE pe24_10(.x(x10),.w(w24_9),.acc(r24_9),.res(r24_10),.clk(clk),.wout(w24_10));
	PE pe24_11(.x(x11),.w(w24_10),.acc(r24_10),.res(r24_11),.clk(clk),.wout(w24_11));
	PE pe24_12(.x(x12),.w(w24_11),.acc(r24_11),.res(r24_12),.clk(clk),.wout(w24_12));
	PE pe24_13(.x(x13),.w(w24_12),.acc(r24_12),.res(r24_13),.clk(clk),.wout(w24_13));
	PE pe24_14(.x(x14),.w(w24_13),.acc(r24_13),.res(r24_14),.clk(clk),.wout(w24_14));
	PE pe24_15(.x(x15),.w(w24_14),.acc(r24_14),.res(r24_15),.clk(clk),.wout(w24_15));
	PE pe24_16(.x(x16),.w(w24_15),.acc(r24_15),.res(r24_16),.clk(clk),.wout(w24_16));
	PE pe24_17(.x(x17),.w(w24_16),.acc(r24_16),.res(r24_17),.clk(clk),.wout(w24_17));
	PE pe24_18(.x(x18),.w(w24_17),.acc(r24_17),.res(r24_18),.clk(clk),.wout(w24_18));
	PE pe24_19(.x(x19),.w(w24_18),.acc(r24_18),.res(r24_19),.clk(clk),.wout(w24_19));
	PE pe24_20(.x(x20),.w(w24_19),.acc(r24_19),.res(r24_20),.clk(clk),.wout(w24_20));
	PE pe24_21(.x(x21),.w(w24_20),.acc(r24_20),.res(r24_21),.clk(clk),.wout(w24_21));
	PE pe24_22(.x(x22),.w(w24_21),.acc(r24_21),.res(r24_22),.clk(clk),.wout(w24_22));
	PE pe24_23(.x(x23),.w(w24_22),.acc(r24_22),.res(r24_23),.clk(clk),.wout(w24_23));
	PE pe24_24(.x(x24),.w(w24_23),.acc(r24_23),.res(r24_24),.clk(clk),.wout(w24_24));
	PE pe24_25(.x(x25),.w(w24_24),.acc(r24_24),.res(r24_25),.clk(clk),.wout(w24_25));
	PE pe24_26(.x(x26),.w(w24_25),.acc(r24_25),.res(r24_26),.clk(clk),.wout(w24_26));
	PE pe24_27(.x(x27),.w(w24_26),.acc(r24_26),.res(r24_27),.clk(clk),.wout(w24_27));
	PE pe24_28(.x(x28),.w(w24_27),.acc(r24_27),.res(r24_28),.clk(clk),.wout(w24_28));
	PE pe24_29(.x(x29),.w(w24_28),.acc(r24_28),.res(r24_29),.clk(clk),.wout(w24_29));
	PE pe24_30(.x(x30),.w(w24_29),.acc(r24_29),.res(r24_30),.clk(clk),.wout(w24_30));
	PE pe24_31(.x(x31),.w(w24_30),.acc(r24_30),.res(r24_31),.clk(clk),.wout(w24_31));
	PE pe24_32(.x(x32),.w(w24_31),.acc(r24_31),.res(r24_32),.clk(clk),.wout(w24_32));
	PE pe24_33(.x(x33),.w(w24_32),.acc(r24_32),.res(r24_33),.clk(clk),.wout(w24_33));
	PE pe24_34(.x(x34),.w(w24_33),.acc(r24_33),.res(r24_34),.clk(clk),.wout(w24_34));
	PE pe24_35(.x(x35),.w(w24_34),.acc(r24_34),.res(r24_35),.clk(clk),.wout(w24_35));
	PE pe24_36(.x(x36),.w(w24_35),.acc(r24_35),.res(r24_36),.clk(clk),.wout(w24_36));
	PE pe24_37(.x(x37),.w(w24_36),.acc(r24_36),.res(r24_37),.clk(clk),.wout(w24_37));
	PE pe24_38(.x(x38),.w(w24_37),.acc(r24_37),.res(r24_38),.clk(clk),.wout(w24_38));
	PE pe24_39(.x(x39),.w(w24_38),.acc(r24_38),.res(r24_39),.clk(clk),.wout(w24_39));
	PE pe24_40(.x(x40),.w(w24_39),.acc(r24_39),.res(r24_40),.clk(clk),.wout(w24_40));
	PE pe24_41(.x(x41),.w(w24_40),.acc(r24_40),.res(r24_41),.clk(clk),.wout(w24_41));
	PE pe24_42(.x(x42),.w(w24_41),.acc(r24_41),.res(r24_42),.clk(clk),.wout(w24_42));
	PE pe24_43(.x(x43),.w(w24_42),.acc(r24_42),.res(r24_43),.clk(clk),.wout(w24_43));
	PE pe24_44(.x(x44),.w(w24_43),.acc(r24_43),.res(r24_44),.clk(clk),.wout(w24_44));
	PE pe24_45(.x(x45),.w(w24_44),.acc(r24_44),.res(r24_45),.clk(clk),.wout(w24_45));
	PE pe24_46(.x(x46),.w(w24_45),.acc(r24_45),.res(r24_46),.clk(clk),.wout(w24_46));
	PE pe24_47(.x(x47),.w(w24_46),.acc(r24_46),.res(r24_47),.clk(clk),.wout(w24_47));
	PE pe24_48(.x(x48),.w(w24_47),.acc(r24_47),.res(r24_48),.clk(clk),.wout(w24_48));
	PE pe24_49(.x(x49),.w(w24_48),.acc(r24_48),.res(r24_49),.clk(clk),.wout(w24_49));
	PE pe24_50(.x(x50),.w(w24_49),.acc(r24_49),.res(r24_50),.clk(clk),.wout(w24_50));
	PE pe24_51(.x(x51),.w(w24_50),.acc(r24_50),.res(r24_51),.clk(clk),.wout(w24_51));
	PE pe24_52(.x(x52),.w(w24_51),.acc(r24_51),.res(r24_52),.clk(clk),.wout(w24_52));
	PE pe24_53(.x(x53),.w(w24_52),.acc(r24_52),.res(r24_53),.clk(clk),.wout(w24_53));
	PE pe24_54(.x(x54),.w(w24_53),.acc(r24_53),.res(r24_54),.clk(clk),.wout(w24_54));
	PE pe24_55(.x(x55),.w(w24_54),.acc(r24_54),.res(r24_55),.clk(clk),.wout(w24_55));
	PE pe24_56(.x(x56),.w(w24_55),.acc(r24_55),.res(r24_56),.clk(clk),.wout(w24_56));
	PE pe24_57(.x(x57),.w(w24_56),.acc(r24_56),.res(r24_57),.clk(clk),.wout(w24_57));
	PE pe24_58(.x(x58),.w(w24_57),.acc(r24_57),.res(r24_58),.clk(clk),.wout(w24_58));
	PE pe24_59(.x(x59),.w(w24_58),.acc(r24_58),.res(r24_59),.clk(clk),.wout(w24_59));
	PE pe24_60(.x(x60),.w(w24_59),.acc(r24_59),.res(r24_60),.clk(clk),.wout(w24_60));
	PE pe24_61(.x(x61),.w(w24_60),.acc(r24_60),.res(r24_61),.clk(clk),.wout(w24_61));
	PE pe24_62(.x(x62),.w(w24_61),.acc(r24_61),.res(r24_62),.clk(clk),.wout(w24_62));
	PE pe24_63(.x(x63),.w(w24_62),.acc(r24_62),.res(r24_63),.clk(clk),.wout(w24_63));
	PE pe24_64(.x(x64),.w(w24_63),.acc(r24_63),.res(r24_64),.clk(clk),.wout(w24_64));
	PE pe24_65(.x(x65),.w(w24_64),.acc(r24_64),.res(r24_65),.clk(clk),.wout(w24_65));
	PE pe24_66(.x(x66),.w(w24_65),.acc(r24_65),.res(r24_66),.clk(clk),.wout(w24_66));
	PE pe24_67(.x(x67),.w(w24_66),.acc(r24_66),.res(r24_67),.clk(clk),.wout(w24_67));
	PE pe24_68(.x(x68),.w(w24_67),.acc(r24_67),.res(r24_68),.clk(clk),.wout(w24_68));
	PE pe24_69(.x(x69),.w(w24_68),.acc(r24_68),.res(r24_69),.clk(clk),.wout(w24_69));
	PE pe24_70(.x(x70),.w(w24_69),.acc(r24_69),.res(r24_70),.clk(clk),.wout(w24_70));
	PE pe24_71(.x(x71),.w(w24_70),.acc(r24_70),.res(r24_71),.clk(clk),.wout(w24_71));
	PE pe24_72(.x(x72),.w(w24_71),.acc(r24_71),.res(r24_72),.clk(clk),.wout(w24_72));
	PE pe24_73(.x(x73),.w(w24_72),.acc(r24_72),.res(r24_73),.clk(clk),.wout(w24_73));
	PE pe24_74(.x(x74),.w(w24_73),.acc(r24_73),.res(r24_74),.clk(clk),.wout(w24_74));
	PE pe24_75(.x(x75),.w(w24_74),.acc(r24_74),.res(r24_75),.clk(clk),.wout(w24_75));
	PE pe24_76(.x(x76),.w(w24_75),.acc(r24_75),.res(r24_76),.clk(clk),.wout(w24_76));
	PE pe24_77(.x(x77),.w(w24_76),.acc(r24_76),.res(r24_77),.clk(clk),.wout(w24_77));
	PE pe24_78(.x(x78),.w(w24_77),.acc(r24_77),.res(r24_78),.clk(clk),.wout(w24_78));
	PE pe24_79(.x(x79),.w(w24_78),.acc(r24_78),.res(r24_79),.clk(clk),.wout(w24_79));
	PE pe24_80(.x(x80),.w(w24_79),.acc(r24_79),.res(r24_80),.clk(clk),.wout(w24_80));
	PE pe24_81(.x(x81),.w(w24_80),.acc(r24_80),.res(r24_81),.clk(clk),.wout(w24_81));
	PE pe24_82(.x(x82),.w(w24_81),.acc(r24_81),.res(r24_82),.clk(clk),.wout(w24_82));
	PE pe24_83(.x(x83),.w(w24_82),.acc(r24_82),.res(r24_83),.clk(clk),.wout(w24_83));
	PE pe24_84(.x(x84),.w(w24_83),.acc(r24_83),.res(r24_84),.clk(clk),.wout(w24_84));
	PE pe24_85(.x(x85),.w(w24_84),.acc(r24_84),.res(r24_85),.clk(clk),.wout(w24_85));
	PE pe24_86(.x(x86),.w(w24_85),.acc(r24_85),.res(r24_86),.clk(clk),.wout(w24_86));
	PE pe24_87(.x(x87),.w(w24_86),.acc(r24_86),.res(r24_87),.clk(clk),.wout(w24_87));
	PE pe24_88(.x(x88),.w(w24_87),.acc(r24_87),.res(r24_88),.clk(clk),.wout(w24_88));
	PE pe24_89(.x(x89),.w(w24_88),.acc(r24_88),.res(r24_89),.clk(clk),.wout(w24_89));
	PE pe24_90(.x(x90),.w(w24_89),.acc(r24_89),.res(r24_90),.clk(clk),.wout(w24_90));
	PE pe24_91(.x(x91),.w(w24_90),.acc(r24_90),.res(r24_91),.clk(clk),.wout(w24_91));
	PE pe24_92(.x(x92),.w(w24_91),.acc(r24_91),.res(r24_92),.clk(clk),.wout(w24_92));
	PE pe24_93(.x(x93),.w(w24_92),.acc(r24_92),.res(r24_93),.clk(clk),.wout(w24_93));
	PE pe24_94(.x(x94),.w(w24_93),.acc(r24_93),.res(r24_94),.clk(clk),.wout(w24_94));
	PE pe24_95(.x(x95),.w(w24_94),.acc(r24_94),.res(r24_95),.clk(clk),.wout(w24_95));
	PE pe24_96(.x(x96),.w(w24_95),.acc(r24_95),.res(r24_96),.clk(clk),.wout(w24_96));
	PE pe24_97(.x(x97),.w(w24_96),.acc(r24_96),.res(r24_97),.clk(clk),.wout(w24_97));
	PE pe24_98(.x(x98),.w(w24_97),.acc(r24_97),.res(r24_98),.clk(clk),.wout(w24_98));
	PE pe24_99(.x(x99),.w(w24_98),.acc(r24_98),.res(r24_99),.clk(clk),.wout(w24_99));
	PE pe24_100(.x(x100),.w(w24_99),.acc(r24_99),.res(r24_100),.clk(clk),.wout(w24_100));
	PE pe24_101(.x(x101),.w(w24_100),.acc(r24_100),.res(r24_101),.clk(clk),.wout(w24_101));
	PE pe24_102(.x(x102),.w(w24_101),.acc(r24_101),.res(r24_102),.clk(clk),.wout(w24_102));
	PE pe24_103(.x(x103),.w(w24_102),.acc(r24_102),.res(r24_103),.clk(clk),.wout(w24_103));
	PE pe24_104(.x(x104),.w(w24_103),.acc(r24_103),.res(r24_104),.clk(clk),.wout(w24_104));
	PE pe24_105(.x(x105),.w(w24_104),.acc(r24_104),.res(r24_105),.clk(clk),.wout(w24_105));
	PE pe24_106(.x(x106),.w(w24_105),.acc(r24_105),.res(r24_106),.clk(clk),.wout(w24_106));
	PE pe24_107(.x(x107),.w(w24_106),.acc(r24_106),.res(r24_107),.clk(clk),.wout(w24_107));
	PE pe24_108(.x(x108),.w(w24_107),.acc(r24_107),.res(r24_108),.clk(clk),.wout(w24_108));
	PE pe24_109(.x(x109),.w(w24_108),.acc(r24_108),.res(r24_109),.clk(clk),.wout(w24_109));
	PE pe24_110(.x(x110),.w(w24_109),.acc(r24_109),.res(r24_110),.clk(clk),.wout(w24_110));
	PE pe24_111(.x(x111),.w(w24_110),.acc(r24_110),.res(r24_111),.clk(clk),.wout(w24_111));
	PE pe24_112(.x(x112),.w(w24_111),.acc(r24_111),.res(r24_112),.clk(clk),.wout(w24_112));
	PE pe24_113(.x(x113),.w(w24_112),.acc(r24_112),.res(r24_113),.clk(clk),.wout(w24_113));
	PE pe24_114(.x(x114),.w(w24_113),.acc(r24_113),.res(r24_114),.clk(clk),.wout(w24_114));
	PE pe24_115(.x(x115),.w(w24_114),.acc(r24_114),.res(r24_115),.clk(clk),.wout(w24_115));
	PE pe24_116(.x(x116),.w(w24_115),.acc(r24_115),.res(r24_116),.clk(clk),.wout(w24_116));
	PE pe24_117(.x(x117),.w(w24_116),.acc(r24_116),.res(r24_117),.clk(clk),.wout(w24_117));
	PE pe24_118(.x(x118),.w(w24_117),.acc(r24_117),.res(r24_118),.clk(clk),.wout(w24_118));
	PE pe24_119(.x(x119),.w(w24_118),.acc(r24_118),.res(r24_119),.clk(clk),.wout(w24_119));
	PE pe24_120(.x(x120),.w(w24_119),.acc(r24_119),.res(r24_120),.clk(clk),.wout(w24_120));
	PE pe24_121(.x(x121),.w(w24_120),.acc(r24_120),.res(r24_121),.clk(clk),.wout(w24_121));
	PE pe24_122(.x(x122),.w(w24_121),.acc(r24_121),.res(r24_122),.clk(clk),.wout(w24_122));
	PE pe24_123(.x(x123),.w(w24_122),.acc(r24_122),.res(r24_123),.clk(clk),.wout(w24_123));
	PE pe24_124(.x(x124),.w(w24_123),.acc(r24_123),.res(r24_124),.clk(clk),.wout(w24_124));
	PE pe24_125(.x(x125),.w(w24_124),.acc(r24_124),.res(r24_125),.clk(clk),.wout(w24_125));
	PE pe24_126(.x(x126),.w(w24_125),.acc(r24_125),.res(r24_126),.clk(clk),.wout(w24_126));
	PE pe24_127(.x(x127),.w(w24_126),.acc(r24_126),.res(result24),.clk(clk),.wout(weight24));

	PE pe25_0(.x(x0),.w(w25),.acc(32'h0),.res(r25_0),.clk(clk),.wout(w25_0));
	PE pe25_1(.x(x1),.w(w25_0),.acc(r25_0),.res(r25_1),.clk(clk),.wout(w25_1));
	PE pe25_2(.x(x2),.w(w25_1),.acc(r25_1),.res(r25_2),.clk(clk),.wout(w25_2));
	PE pe25_3(.x(x3),.w(w25_2),.acc(r25_2),.res(r25_3),.clk(clk),.wout(w25_3));
	PE pe25_4(.x(x4),.w(w25_3),.acc(r25_3),.res(r25_4),.clk(clk),.wout(w25_4));
	PE pe25_5(.x(x5),.w(w25_4),.acc(r25_4),.res(r25_5),.clk(clk),.wout(w25_5));
	PE pe25_6(.x(x6),.w(w25_5),.acc(r25_5),.res(r25_6),.clk(clk),.wout(w25_6));
	PE pe25_7(.x(x7),.w(w25_6),.acc(r25_6),.res(r25_7),.clk(clk),.wout(w25_7));
	PE pe25_8(.x(x8),.w(w25_7),.acc(r25_7),.res(r25_8),.clk(clk),.wout(w25_8));
	PE pe25_9(.x(x9),.w(w25_8),.acc(r25_8),.res(r25_9),.clk(clk),.wout(w25_9));
	PE pe25_10(.x(x10),.w(w25_9),.acc(r25_9),.res(r25_10),.clk(clk),.wout(w25_10));
	PE pe25_11(.x(x11),.w(w25_10),.acc(r25_10),.res(r25_11),.clk(clk),.wout(w25_11));
	PE pe25_12(.x(x12),.w(w25_11),.acc(r25_11),.res(r25_12),.clk(clk),.wout(w25_12));
	PE pe25_13(.x(x13),.w(w25_12),.acc(r25_12),.res(r25_13),.clk(clk),.wout(w25_13));
	PE pe25_14(.x(x14),.w(w25_13),.acc(r25_13),.res(r25_14),.clk(clk),.wout(w25_14));
	PE pe25_15(.x(x15),.w(w25_14),.acc(r25_14),.res(r25_15),.clk(clk),.wout(w25_15));
	PE pe25_16(.x(x16),.w(w25_15),.acc(r25_15),.res(r25_16),.clk(clk),.wout(w25_16));
	PE pe25_17(.x(x17),.w(w25_16),.acc(r25_16),.res(r25_17),.clk(clk),.wout(w25_17));
	PE pe25_18(.x(x18),.w(w25_17),.acc(r25_17),.res(r25_18),.clk(clk),.wout(w25_18));
	PE pe25_19(.x(x19),.w(w25_18),.acc(r25_18),.res(r25_19),.clk(clk),.wout(w25_19));
	PE pe25_20(.x(x20),.w(w25_19),.acc(r25_19),.res(r25_20),.clk(clk),.wout(w25_20));
	PE pe25_21(.x(x21),.w(w25_20),.acc(r25_20),.res(r25_21),.clk(clk),.wout(w25_21));
	PE pe25_22(.x(x22),.w(w25_21),.acc(r25_21),.res(r25_22),.clk(clk),.wout(w25_22));
	PE pe25_23(.x(x23),.w(w25_22),.acc(r25_22),.res(r25_23),.clk(clk),.wout(w25_23));
	PE pe25_24(.x(x24),.w(w25_23),.acc(r25_23),.res(r25_24),.clk(clk),.wout(w25_24));
	PE pe25_25(.x(x25),.w(w25_24),.acc(r25_24),.res(r25_25),.clk(clk),.wout(w25_25));
	PE pe25_26(.x(x26),.w(w25_25),.acc(r25_25),.res(r25_26),.clk(clk),.wout(w25_26));
	PE pe25_27(.x(x27),.w(w25_26),.acc(r25_26),.res(r25_27),.clk(clk),.wout(w25_27));
	PE pe25_28(.x(x28),.w(w25_27),.acc(r25_27),.res(r25_28),.clk(clk),.wout(w25_28));
	PE pe25_29(.x(x29),.w(w25_28),.acc(r25_28),.res(r25_29),.clk(clk),.wout(w25_29));
	PE pe25_30(.x(x30),.w(w25_29),.acc(r25_29),.res(r25_30),.clk(clk),.wout(w25_30));
	PE pe25_31(.x(x31),.w(w25_30),.acc(r25_30),.res(r25_31),.clk(clk),.wout(w25_31));
	PE pe25_32(.x(x32),.w(w25_31),.acc(r25_31),.res(r25_32),.clk(clk),.wout(w25_32));
	PE pe25_33(.x(x33),.w(w25_32),.acc(r25_32),.res(r25_33),.clk(clk),.wout(w25_33));
	PE pe25_34(.x(x34),.w(w25_33),.acc(r25_33),.res(r25_34),.clk(clk),.wout(w25_34));
	PE pe25_35(.x(x35),.w(w25_34),.acc(r25_34),.res(r25_35),.clk(clk),.wout(w25_35));
	PE pe25_36(.x(x36),.w(w25_35),.acc(r25_35),.res(r25_36),.clk(clk),.wout(w25_36));
	PE pe25_37(.x(x37),.w(w25_36),.acc(r25_36),.res(r25_37),.clk(clk),.wout(w25_37));
	PE pe25_38(.x(x38),.w(w25_37),.acc(r25_37),.res(r25_38),.clk(clk),.wout(w25_38));
	PE pe25_39(.x(x39),.w(w25_38),.acc(r25_38),.res(r25_39),.clk(clk),.wout(w25_39));
	PE pe25_40(.x(x40),.w(w25_39),.acc(r25_39),.res(r25_40),.clk(clk),.wout(w25_40));
	PE pe25_41(.x(x41),.w(w25_40),.acc(r25_40),.res(r25_41),.clk(clk),.wout(w25_41));
	PE pe25_42(.x(x42),.w(w25_41),.acc(r25_41),.res(r25_42),.clk(clk),.wout(w25_42));
	PE pe25_43(.x(x43),.w(w25_42),.acc(r25_42),.res(r25_43),.clk(clk),.wout(w25_43));
	PE pe25_44(.x(x44),.w(w25_43),.acc(r25_43),.res(r25_44),.clk(clk),.wout(w25_44));
	PE pe25_45(.x(x45),.w(w25_44),.acc(r25_44),.res(r25_45),.clk(clk),.wout(w25_45));
	PE pe25_46(.x(x46),.w(w25_45),.acc(r25_45),.res(r25_46),.clk(clk),.wout(w25_46));
	PE pe25_47(.x(x47),.w(w25_46),.acc(r25_46),.res(r25_47),.clk(clk),.wout(w25_47));
	PE pe25_48(.x(x48),.w(w25_47),.acc(r25_47),.res(r25_48),.clk(clk),.wout(w25_48));
	PE pe25_49(.x(x49),.w(w25_48),.acc(r25_48),.res(r25_49),.clk(clk),.wout(w25_49));
	PE pe25_50(.x(x50),.w(w25_49),.acc(r25_49),.res(r25_50),.clk(clk),.wout(w25_50));
	PE pe25_51(.x(x51),.w(w25_50),.acc(r25_50),.res(r25_51),.clk(clk),.wout(w25_51));
	PE pe25_52(.x(x52),.w(w25_51),.acc(r25_51),.res(r25_52),.clk(clk),.wout(w25_52));
	PE pe25_53(.x(x53),.w(w25_52),.acc(r25_52),.res(r25_53),.clk(clk),.wout(w25_53));
	PE pe25_54(.x(x54),.w(w25_53),.acc(r25_53),.res(r25_54),.clk(clk),.wout(w25_54));
	PE pe25_55(.x(x55),.w(w25_54),.acc(r25_54),.res(r25_55),.clk(clk),.wout(w25_55));
	PE pe25_56(.x(x56),.w(w25_55),.acc(r25_55),.res(r25_56),.clk(clk),.wout(w25_56));
	PE pe25_57(.x(x57),.w(w25_56),.acc(r25_56),.res(r25_57),.clk(clk),.wout(w25_57));
	PE pe25_58(.x(x58),.w(w25_57),.acc(r25_57),.res(r25_58),.clk(clk),.wout(w25_58));
	PE pe25_59(.x(x59),.w(w25_58),.acc(r25_58),.res(r25_59),.clk(clk),.wout(w25_59));
	PE pe25_60(.x(x60),.w(w25_59),.acc(r25_59),.res(r25_60),.clk(clk),.wout(w25_60));
	PE pe25_61(.x(x61),.w(w25_60),.acc(r25_60),.res(r25_61),.clk(clk),.wout(w25_61));
	PE pe25_62(.x(x62),.w(w25_61),.acc(r25_61),.res(r25_62),.clk(clk),.wout(w25_62));
	PE pe25_63(.x(x63),.w(w25_62),.acc(r25_62),.res(r25_63),.clk(clk),.wout(w25_63));
	PE pe25_64(.x(x64),.w(w25_63),.acc(r25_63),.res(r25_64),.clk(clk),.wout(w25_64));
	PE pe25_65(.x(x65),.w(w25_64),.acc(r25_64),.res(r25_65),.clk(clk),.wout(w25_65));
	PE pe25_66(.x(x66),.w(w25_65),.acc(r25_65),.res(r25_66),.clk(clk),.wout(w25_66));
	PE pe25_67(.x(x67),.w(w25_66),.acc(r25_66),.res(r25_67),.clk(clk),.wout(w25_67));
	PE pe25_68(.x(x68),.w(w25_67),.acc(r25_67),.res(r25_68),.clk(clk),.wout(w25_68));
	PE pe25_69(.x(x69),.w(w25_68),.acc(r25_68),.res(r25_69),.clk(clk),.wout(w25_69));
	PE pe25_70(.x(x70),.w(w25_69),.acc(r25_69),.res(r25_70),.clk(clk),.wout(w25_70));
	PE pe25_71(.x(x71),.w(w25_70),.acc(r25_70),.res(r25_71),.clk(clk),.wout(w25_71));
	PE pe25_72(.x(x72),.w(w25_71),.acc(r25_71),.res(r25_72),.clk(clk),.wout(w25_72));
	PE pe25_73(.x(x73),.w(w25_72),.acc(r25_72),.res(r25_73),.clk(clk),.wout(w25_73));
	PE pe25_74(.x(x74),.w(w25_73),.acc(r25_73),.res(r25_74),.clk(clk),.wout(w25_74));
	PE pe25_75(.x(x75),.w(w25_74),.acc(r25_74),.res(r25_75),.clk(clk),.wout(w25_75));
	PE pe25_76(.x(x76),.w(w25_75),.acc(r25_75),.res(r25_76),.clk(clk),.wout(w25_76));
	PE pe25_77(.x(x77),.w(w25_76),.acc(r25_76),.res(r25_77),.clk(clk),.wout(w25_77));
	PE pe25_78(.x(x78),.w(w25_77),.acc(r25_77),.res(r25_78),.clk(clk),.wout(w25_78));
	PE pe25_79(.x(x79),.w(w25_78),.acc(r25_78),.res(r25_79),.clk(clk),.wout(w25_79));
	PE pe25_80(.x(x80),.w(w25_79),.acc(r25_79),.res(r25_80),.clk(clk),.wout(w25_80));
	PE pe25_81(.x(x81),.w(w25_80),.acc(r25_80),.res(r25_81),.clk(clk),.wout(w25_81));
	PE pe25_82(.x(x82),.w(w25_81),.acc(r25_81),.res(r25_82),.clk(clk),.wout(w25_82));
	PE pe25_83(.x(x83),.w(w25_82),.acc(r25_82),.res(r25_83),.clk(clk),.wout(w25_83));
	PE pe25_84(.x(x84),.w(w25_83),.acc(r25_83),.res(r25_84),.clk(clk),.wout(w25_84));
	PE pe25_85(.x(x85),.w(w25_84),.acc(r25_84),.res(r25_85),.clk(clk),.wout(w25_85));
	PE pe25_86(.x(x86),.w(w25_85),.acc(r25_85),.res(r25_86),.clk(clk),.wout(w25_86));
	PE pe25_87(.x(x87),.w(w25_86),.acc(r25_86),.res(r25_87),.clk(clk),.wout(w25_87));
	PE pe25_88(.x(x88),.w(w25_87),.acc(r25_87),.res(r25_88),.clk(clk),.wout(w25_88));
	PE pe25_89(.x(x89),.w(w25_88),.acc(r25_88),.res(r25_89),.clk(clk),.wout(w25_89));
	PE pe25_90(.x(x90),.w(w25_89),.acc(r25_89),.res(r25_90),.clk(clk),.wout(w25_90));
	PE pe25_91(.x(x91),.w(w25_90),.acc(r25_90),.res(r25_91),.clk(clk),.wout(w25_91));
	PE pe25_92(.x(x92),.w(w25_91),.acc(r25_91),.res(r25_92),.clk(clk),.wout(w25_92));
	PE pe25_93(.x(x93),.w(w25_92),.acc(r25_92),.res(r25_93),.clk(clk),.wout(w25_93));
	PE pe25_94(.x(x94),.w(w25_93),.acc(r25_93),.res(r25_94),.clk(clk),.wout(w25_94));
	PE pe25_95(.x(x95),.w(w25_94),.acc(r25_94),.res(r25_95),.clk(clk),.wout(w25_95));
	PE pe25_96(.x(x96),.w(w25_95),.acc(r25_95),.res(r25_96),.clk(clk),.wout(w25_96));
	PE pe25_97(.x(x97),.w(w25_96),.acc(r25_96),.res(r25_97),.clk(clk),.wout(w25_97));
	PE pe25_98(.x(x98),.w(w25_97),.acc(r25_97),.res(r25_98),.clk(clk),.wout(w25_98));
	PE pe25_99(.x(x99),.w(w25_98),.acc(r25_98),.res(r25_99),.clk(clk),.wout(w25_99));
	PE pe25_100(.x(x100),.w(w25_99),.acc(r25_99),.res(r25_100),.clk(clk),.wout(w25_100));
	PE pe25_101(.x(x101),.w(w25_100),.acc(r25_100),.res(r25_101),.clk(clk),.wout(w25_101));
	PE pe25_102(.x(x102),.w(w25_101),.acc(r25_101),.res(r25_102),.clk(clk),.wout(w25_102));
	PE pe25_103(.x(x103),.w(w25_102),.acc(r25_102),.res(r25_103),.clk(clk),.wout(w25_103));
	PE pe25_104(.x(x104),.w(w25_103),.acc(r25_103),.res(r25_104),.clk(clk),.wout(w25_104));
	PE pe25_105(.x(x105),.w(w25_104),.acc(r25_104),.res(r25_105),.clk(clk),.wout(w25_105));
	PE pe25_106(.x(x106),.w(w25_105),.acc(r25_105),.res(r25_106),.clk(clk),.wout(w25_106));
	PE pe25_107(.x(x107),.w(w25_106),.acc(r25_106),.res(r25_107),.clk(clk),.wout(w25_107));
	PE pe25_108(.x(x108),.w(w25_107),.acc(r25_107),.res(r25_108),.clk(clk),.wout(w25_108));
	PE pe25_109(.x(x109),.w(w25_108),.acc(r25_108),.res(r25_109),.clk(clk),.wout(w25_109));
	PE pe25_110(.x(x110),.w(w25_109),.acc(r25_109),.res(r25_110),.clk(clk),.wout(w25_110));
	PE pe25_111(.x(x111),.w(w25_110),.acc(r25_110),.res(r25_111),.clk(clk),.wout(w25_111));
	PE pe25_112(.x(x112),.w(w25_111),.acc(r25_111),.res(r25_112),.clk(clk),.wout(w25_112));
	PE pe25_113(.x(x113),.w(w25_112),.acc(r25_112),.res(r25_113),.clk(clk),.wout(w25_113));
	PE pe25_114(.x(x114),.w(w25_113),.acc(r25_113),.res(r25_114),.clk(clk),.wout(w25_114));
	PE pe25_115(.x(x115),.w(w25_114),.acc(r25_114),.res(r25_115),.clk(clk),.wout(w25_115));
	PE pe25_116(.x(x116),.w(w25_115),.acc(r25_115),.res(r25_116),.clk(clk),.wout(w25_116));
	PE pe25_117(.x(x117),.w(w25_116),.acc(r25_116),.res(r25_117),.clk(clk),.wout(w25_117));
	PE pe25_118(.x(x118),.w(w25_117),.acc(r25_117),.res(r25_118),.clk(clk),.wout(w25_118));
	PE pe25_119(.x(x119),.w(w25_118),.acc(r25_118),.res(r25_119),.clk(clk),.wout(w25_119));
	PE pe25_120(.x(x120),.w(w25_119),.acc(r25_119),.res(r25_120),.clk(clk),.wout(w25_120));
	PE pe25_121(.x(x121),.w(w25_120),.acc(r25_120),.res(r25_121),.clk(clk),.wout(w25_121));
	PE pe25_122(.x(x122),.w(w25_121),.acc(r25_121),.res(r25_122),.clk(clk),.wout(w25_122));
	PE pe25_123(.x(x123),.w(w25_122),.acc(r25_122),.res(r25_123),.clk(clk),.wout(w25_123));
	PE pe25_124(.x(x124),.w(w25_123),.acc(r25_123),.res(r25_124),.clk(clk),.wout(w25_124));
	PE pe25_125(.x(x125),.w(w25_124),.acc(r25_124),.res(r25_125),.clk(clk),.wout(w25_125));
	PE pe25_126(.x(x126),.w(w25_125),.acc(r25_125),.res(r25_126),.clk(clk),.wout(w25_126));
	PE pe25_127(.x(x127),.w(w25_126),.acc(r25_126),.res(result25),.clk(clk),.wout(weight25));

	PE pe26_0(.x(x0),.w(w26),.acc(32'h0),.res(r26_0),.clk(clk),.wout(w26_0));
	PE pe26_1(.x(x1),.w(w26_0),.acc(r26_0),.res(r26_1),.clk(clk),.wout(w26_1));
	PE pe26_2(.x(x2),.w(w26_1),.acc(r26_1),.res(r26_2),.clk(clk),.wout(w26_2));
	PE pe26_3(.x(x3),.w(w26_2),.acc(r26_2),.res(r26_3),.clk(clk),.wout(w26_3));
	PE pe26_4(.x(x4),.w(w26_3),.acc(r26_3),.res(r26_4),.clk(clk),.wout(w26_4));
	PE pe26_5(.x(x5),.w(w26_4),.acc(r26_4),.res(r26_5),.clk(clk),.wout(w26_5));
	PE pe26_6(.x(x6),.w(w26_5),.acc(r26_5),.res(r26_6),.clk(clk),.wout(w26_6));
	PE pe26_7(.x(x7),.w(w26_6),.acc(r26_6),.res(r26_7),.clk(clk),.wout(w26_7));
	PE pe26_8(.x(x8),.w(w26_7),.acc(r26_7),.res(r26_8),.clk(clk),.wout(w26_8));
	PE pe26_9(.x(x9),.w(w26_8),.acc(r26_8),.res(r26_9),.clk(clk),.wout(w26_9));
	PE pe26_10(.x(x10),.w(w26_9),.acc(r26_9),.res(r26_10),.clk(clk),.wout(w26_10));
	PE pe26_11(.x(x11),.w(w26_10),.acc(r26_10),.res(r26_11),.clk(clk),.wout(w26_11));
	PE pe26_12(.x(x12),.w(w26_11),.acc(r26_11),.res(r26_12),.clk(clk),.wout(w26_12));
	PE pe26_13(.x(x13),.w(w26_12),.acc(r26_12),.res(r26_13),.clk(clk),.wout(w26_13));
	PE pe26_14(.x(x14),.w(w26_13),.acc(r26_13),.res(r26_14),.clk(clk),.wout(w26_14));
	PE pe26_15(.x(x15),.w(w26_14),.acc(r26_14),.res(r26_15),.clk(clk),.wout(w26_15));
	PE pe26_16(.x(x16),.w(w26_15),.acc(r26_15),.res(r26_16),.clk(clk),.wout(w26_16));
	PE pe26_17(.x(x17),.w(w26_16),.acc(r26_16),.res(r26_17),.clk(clk),.wout(w26_17));
	PE pe26_18(.x(x18),.w(w26_17),.acc(r26_17),.res(r26_18),.clk(clk),.wout(w26_18));
	PE pe26_19(.x(x19),.w(w26_18),.acc(r26_18),.res(r26_19),.clk(clk),.wout(w26_19));
	PE pe26_20(.x(x20),.w(w26_19),.acc(r26_19),.res(r26_20),.clk(clk),.wout(w26_20));
	PE pe26_21(.x(x21),.w(w26_20),.acc(r26_20),.res(r26_21),.clk(clk),.wout(w26_21));
	PE pe26_22(.x(x22),.w(w26_21),.acc(r26_21),.res(r26_22),.clk(clk),.wout(w26_22));
	PE pe26_23(.x(x23),.w(w26_22),.acc(r26_22),.res(r26_23),.clk(clk),.wout(w26_23));
	PE pe26_24(.x(x24),.w(w26_23),.acc(r26_23),.res(r26_24),.clk(clk),.wout(w26_24));
	PE pe26_25(.x(x25),.w(w26_24),.acc(r26_24),.res(r26_25),.clk(clk),.wout(w26_25));
	PE pe26_26(.x(x26),.w(w26_25),.acc(r26_25),.res(r26_26),.clk(clk),.wout(w26_26));
	PE pe26_27(.x(x27),.w(w26_26),.acc(r26_26),.res(r26_27),.clk(clk),.wout(w26_27));
	PE pe26_28(.x(x28),.w(w26_27),.acc(r26_27),.res(r26_28),.clk(clk),.wout(w26_28));
	PE pe26_29(.x(x29),.w(w26_28),.acc(r26_28),.res(r26_29),.clk(clk),.wout(w26_29));
	PE pe26_30(.x(x30),.w(w26_29),.acc(r26_29),.res(r26_30),.clk(clk),.wout(w26_30));
	PE pe26_31(.x(x31),.w(w26_30),.acc(r26_30),.res(r26_31),.clk(clk),.wout(w26_31));
	PE pe26_32(.x(x32),.w(w26_31),.acc(r26_31),.res(r26_32),.clk(clk),.wout(w26_32));
	PE pe26_33(.x(x33),.w(w26_32),.acc(r26_32),.res(r26_33),.clk(clk),.wout(w26_33));
	PE pe26_34(.x(x34),.w(w26_33),.acc(r26_33),.res(r26_34),.clk(clk),.wout(w26_34));
	PE pe26_35(.x(x35),.w(w26_34),.acc(r26_34),.res(r26_35),.clk(clk),.wout(w26_35));
	PE pe26_36(.x(x36),.w(w26_35),.acc(r26_35),.res(r26_36),.clk(clk),.wout(w26_36));
	PE pe26_37(.x(x37),.w(w26_36),.acc(r26_36),.res(r26_37),.clk(clk),.wout(w26_37));
	PE pe26_38(.x(x38),.w(w26_37),.acc(r26_37),.res(r26_38),.clk(clk),.wout(w26_38));
	PE pe26_39(.x(x39),.w(w26_38),.acc(r26_38),.res(r26_39),.clk(clk),.wout(w26_39));
	PE pe26_40(.x(x40),.w(w26_39),.acc(r26_39),.res(r26_40),.clk(clk),.wout(w26_40));
	PE pe26_41(.x(x41),.w(w26_40),.acc(r26_40),.res(r26_41),.clk(clk),.wout(w26_41));
	PE pe26_42(.x(x42),.w(w26_41),.acc(r26_41),.res(r26_42),.clk(clk),.wout(w26_42));
	PE pe26_43(.x(x43),.w(w26_42),.acc(r26_42),.res(r26_43),.clk(clk),.wout(w26_43));
	PE pe26_44(.x(x44),.w(w26_43),.acc(r26_43),.res(r26_44),.clk(clk),.wout(w26_44));
	PE pe26_45(.x(x45),.w(w26_44),.acc(r26_44),.res(r26_45),.clk(clk),.wout(w26_45));
	PE pe26_46(.x(x46),.w(w26_45),.acc(r26_45),.res(r26_46),.clk(clk),.wout(w26_46));
	PE pe26_47(.x(x47),.w(w26_46),.acc(r26_46),.res(r26_47),.clk(clk),.wout(w26_47));
	PE pe26_48(.x(x48),.w(w26_47),.acc(r26_47),.res(r26_48),.clk(clk),.wout(w26_48));
	PE pe26_49(.x(x49),.w(w26_48),.acc(r26_48),.res(r26_49),.clk(clk),.wout(w26_49));
	PE pe26_50(.x(x50),.w(w26_49),.acc(r26_49),.res(r26_50),.clk(clk),.wout(w26_50));
	PE pe26_51(.x(x51),.w(w26_50),.acc(r26_50),.res(r26_51),.clk(clk),.wout(w26_51));
	PE pe26_52(.x(x52),.w(w26_51),.acc(r26_51),.res(r26_52),.clk(clk),.wout(w26_52));
	PE pe26_53(.x(x53),.w(w26_52),.acc(r26_52),.res(r26_53),.clk(clk),.wout(w26_53));
	PE pe26_54(.x(x54),.w(w26_53),.acc(r26_53),.res(r26_54),.clk(clk),.wout(w26_54));
	PE pe26_55(.x(x55),.w(w26_54),.acc(r26_54),.res(r26_55),.clk(clk),.wout(w26_55));
	PE pe26_56(.x(x56),.w(w26_55),.acc(r26_55),.res(r26_56),.clk(clk),.wout(w26_56));
	PE pe26_57(.x(x57),.w(w26_56),.acc(r26_56),.res(r26_57),.clk(clk),.wout(w26_57));
	PE pe26_58(.x(x58),.w(w26_57),.acc(r26_57),.res(r26_58),.clk(clk),.wout(w26_58));
	PE pe26_59(.x(x59),.w(w26_58),.acc(r26_58),.res(r26_59),.clk(clk),.wout(w26_59));
	PE pe26_60(.x(x60),.w(w26_59),.acc(r26_59),.res(r26_60),.clk(clk),.wout(w26_60));
	PE pe26_61(.x(x61),.w(w26_60),.acc(r26_60),.res(r26_61),.clk(clk),.wout(w26_61));
	PE pe26_62(.x(x62),.w(w26_61),.acc(r26_61),.res(r26_62),.clk(clk),.wout(w26_62));
	PE pe26_63(.x(x63),.w(w26_62),.acc(r26_62),.res(r26_63),.clk(clk),.wout(w26_63));
	PE pe26_64(.x(x64),.w(w26_63),.acc(r26_63),.res(r26_64),.clk(clk),.wout(w26_64));
	PE pe26_65(.x(x65),.w(w26_64),.acc(r26_64),.res(r26_65),.clk(clk),.wout(w26_65));
	PE pe26_66(.x(x66),.w(w26_65),.acc(r26_65),.res(r26_66),.clk(clk),.wout(w26_66));
	PE pe26_67(.x(x67),.w(w26_66),.acc(r26_66),.res(r26_67),.clk(clk),.wout(w26_67));
	PE pe26_68(.x(x68),.w(w26_67),.acc(r26_67),.res(r26_68),.clk(clk),.wout(w26_68));
	PE pe26_69(.x(x69),.w(w26_68),.acc(r26_68),.res(r26_69),.clk(clk),.wout(w26_69));
	PE pe26_70(.x(x70),.w(w26_69),.acc(r26_69),.res(r26_70),.clk(clk),.wout(w26_70));
	PE pe26_71(.x(x71),.w(w26_70),.acc(r26_70),.res(r26_71),.clk(clk),.wout(w26_71));
	PE pe26_72(.x(x72),.w(w26_71),.acc(r26_71),.res(r26_72),.clk(clk),.wout(w26_72));
	PE pe26_73(.x(x73),.w(w26_72),.acc(r26_72),.res(r26_73),.clk(clk),.wout(w26_73));
	PE pe26_74(.x(x74),.w(w26_73),.acc(r26_73),.res(r26_74),.clk(clk),.wout(w26_74));
	PE pe26_75(.x(x75),.w(w26_74),.acc(r26_74),.res(r26_75),.clk(clk),.wout(w26_75));
	PE pe26_76(.x(x76),.w(w26_75),.acc(r26_75),.res(r26_76),.clk(clk),.wout(w26_76));
	PE pe26_77(.x(x77),.w(w26_76),.acc(r26_76),.res(r26_77),.clk(clk),.wout(w26_77));
	PE pe26_78(.x(x78),.w(w26_77),.acc(r26_77),.res(r26_78),.clk(clk),.wout(w26_78));
	PE pe26_79(.x(x79),.w(w26_78),.acc(r26_78),.res(r26_79),.clk(clk),.wout(w26_79));
	PE pe26_80(.x(x80),.w(w26_79),.acc(r26_79),.res(r26_80),.clk(clk),.wout(w26_80));
	PE pe26_81(.x(x81),.w(w26_80),.acc(r26_80),.res(r26_81),.clk(clk),.wout(w26_81));
	PE pe26_82(.x(x82),.w(w26_81),.acc(r26_81),.res(r26_82),.clk(clk),.wout(w26_82));
	PE pe26_83(.x(x83),.w(w26_82),.acc(r26_82),.res(r26_83),.clk(clk),.wout(w26_83));
	PE pe26_84(.x(x84),.w(w26_83),.acc(r26_83),.res(r26_84),.clk(clk),.wout(w26_84));
	PE pe26_85(.x(x85),.w(w26_84),.acc(r26_84),.res(r26_85),.clk(clk),.wout(w26_85));
	PE pe26_86(.x(x86),.w(w26_85),.acc(r26_85),.res(r26_86),.clk(clk),.wout(w26_86));
	PE pe26_87(.x(x87),.w(w26_86),.acc(r26_86),.res(r26_87),.clk(clk),.wout(w26_87));
	PE pe26_88(.x(x88),.w(w26_87),.acc(r26_87),.res(r26_88),.clk(clk),.wout(w26_88));
	PE pe26_89(.x(x89),.w(w26_88),.acc(r26_88),.res(r26_89),.clk(clk),.wout(w26_89));
	PE pe26_90(.x(x90),.w(w26_89),.acc(r26_89),.res(r26_90),.clk(clk),.wout(w26_90));
	PE pe26_91(.x(x91),.w(w26_90),.acc(r26_90),.res(r26_91),.clk(clk),.wout(w26_91));
	PE pe26_92(.x(x92),.w(w26_91),.acc(r26_91),.res(r26_92),.clk(clk),.wout(w26_92));
	PE pe26_93(.x(x93),.w(w26_92),.acc(r26_92),.res(r26_93),.clk(clk),.wout(w26_93));
	PE pe26_94(.x(x94),.w(w26_93),.acc(r26_93),.res(r26_94),.clk(clk),.wout(w26_94));
	PE pe26_95(.x(x95),.w(w26_94),.acc(r26_94),.res(r26_95),.clk(clk),.wout(w26_95));
	PE pe26_96(.x(x96),.w(w26_95),.acc(r26_95),.res(r26_96),.clk(clk),.wout(w26_96));
	PE pe26_97(.x(x97),.w(w26_96),.acc(r26_96),.res(r26_97),.clk(clk),.wout(w26_97));
	PE pe26_98(.x(x98),.w(w26_97),.acc(r26_97),.res(r26_98),.clk(clk),.wout(w26_98));
	PE pe26_99(.x(x99),.w(w26_98),.acc(r26_98),.res(r26_99),.clk(clk),.wout(w26_99));
	PE pe26_100(.x(x100),.w(w26_99),.acc(r26_99),.res(r26_100),.clk(clk),.wout(w26_100));
	PE pe26_101(.x(x101),.w(w26_100),.acc(r26_100),.res(r26_101),.clk(clk),.wout(w26_101));
	PE pe26_102(.x(x102),.w(w26_101),.acc(r26_101),.res(r26_102),.clk(clk),.wout(w26_102));
	PE pe26_103(.x(x103),.w(w26_102),.acc(r26_102),.res(r26_103),.clk(clk),.wout(w26_103));
	PE pe26_104(.x(x104),.w(w26_103),.acc(r26_103),.res(r26_104),.clk(clk),.wout(w26_104));
	PE pe26_105(.x(x105),.w(w26_104),.acc(r26_104),.res(r26_105),.clk(clk),.wout(w26_105));
	PE pe26_106(.x(x106),.w(w26_105),.acc(r26_105),.res(r26_106),.clk(clk),.wout(w26_106));
	PE pe26_107(.x(x107),.w(w26_106),.acc(r26_106),.res(r26_107),.clk(clk),.wout(w26_107));
	PE pe26_108(.x(x108),.w(w26_107),.acc(r26_107),.res(r26_108),.clk(clk),.wout(w26_108));
	PE pe26_109(.x(x109),.w(w26_108),.acc(r26_108),.res(r26_109),.clk(clk),.wout(w26_109));
	PE pe26_110(.x(x110),.w(w26_109),.acc(r26_109),.res(r26_110),.clk(clk),.wout(w26_110));
	PE pe26_111(.x(x111),.w(w26_110),.acc(r26_110),.res(r26_111),.clk(clk),.wout(w26_111));
	PE pe26_112(.x(x112),.w(w26_111),.acc(r26_111),.res(r26_112),.clk(clk),.wout(w26_112));
	PE pe26_113(.x(x113),.w(w26_112),.acc(r26_112),.res(r26_113),.clk(clk),.wout(w26_113));
	PE pe26_114(.x(x114),.w(w26_113),.acc(r26_113),.res(r26_114),.clk(clk),.wout(w26_114));
	PE pe26_115(.x(x115),.w(w26_114),.acc(r26_114),.res(r26_115),.clk(clk),.wout(w26_115));
	PE pe26_116(.x(x116),.w(w26_115),.acc(r26_115),.res(r26_116),.clk(clk),.wout(w26_116));
	PE pe26_117(.x(x117),.w(w26_116),.acc(r26_116),.res(r26_117),.clk(clk),.wout(w26_117));
	PE pe26_118(.x(x118),.w(w26_117),.acc(r26_117),.res(r26_118),.clk(clk),.wout(w26_118));
	PE pe26_119(.x(x119),.w(w26_118),.acc(r26_118),.res(r26_119),.clk(clk),.wout(w26_119));
	PE pe26_120(.x(x120),.w(w26_119),.acc(r26_119),.res(r26_120),.clk(clk),.wout(w26_120));
	PE pe26_121(.x(x121),.w(w26_120),.acc(r26_120),.res(r26_121),.clk(clk),.wout(w26_121));
	PE pe26_122(.x(x122),.w(w26_121),.acc(r26_121),.res(r26_122),.clk(clk),.wout(w26_122));
	PE pe26_123(.x(x123),.w(w26_122),.acc(r26_122),.res(r26_123),.clk(clk),.wout(w26_123));
	PE pe26_124(.x(x124),.w(w26_123),.acc(r26_123),.res(r26_124),.clk(clk),.wout(w26_124));
	PE pe26_125(.x(x125),.w(w26_124),.acc(r26_124),.res(r26_125),.clk(clk),.wout(w26_125));
	PE pe26_126(.x(x126),.w(w26_125),.acc(r26_125),.res(r26_126),.clk(clk),.wout(w26_126));
	PE pe26_127(.x(x127),.w(w26_126),.acc(r26_126),.res(result26),.clk(clk),.wout(weight26));

	PE pe27_0(.x(x0),.w(w27),.acc(32'h0),.res(r27_0),.clk(clk),.wout(w27_0));
	PE pe27_1(.x(x1),.w(w27_0),.acc(r27_0),.res(r27_1),.clk(clk),.wout(w27_1));
	PE pe27_2(.x(x2),.w(w27_1),.acc(r27_1),.res(r27_2),.clk(clk),.wout(w27_2));
	PE pe27_3(.x(x3),.w(w27_2),.acc(r27_2),.res(r27_3),.clk(clk),.wout(w27_3));
	PE pe27_4(.x(x4),.w(w27_3),.acc(r27_3),.res(r27_4),.clk(clk),.wout(w27_4));
	PE pe27_5(.x(x5),.w(w27_4),.acc(r27_4),.res(r27_5),.clk(clk),.wout(w27_5));
	PE pe27_6(.x(x6),.w(w27_5),.acc(r27_5),.res(r27_6),.clk(clk),.wout(w27_6));
	PE pe27_7(.x(x7),.w(w27_6),.acc(r27_6),.res(r27_7),.clk(clk),.wout(w27_7));
	PE pe27_8(.x(x8),.w(w27_7),.acc(r27_7),.res(r27_8),.clk(clk),.wout(w27_8));
	PE pe27_9(.x(x9),.w(w27_8),.acc(r27_8),.res(r27_9),.clk(clk),.wout(w27_9));
	PE pe27_10(.x(x10),.w(w27_9),.acc(r27_9),.res(r27_10),.clk(clk),.wout(w27_10));
	PE pe27_11(.x(x11),.w(w27_10),.acc(r27_10),.res(r27_11),.clk(clk),.wout(w27_11));
	PE pe27_12(.x(x12),.w(w27_11),.acc(r27_11),.res(r27_12),.clk(clk),.wout(w27_12));
	PE pe27_13(.x(x13),.w(w27_12),.acc(r27_12),.res(r27_13),.clk(clk),.wout(w27_13));
	PE pe27_14(.x(x14),.w(w27_13),.acc(r27_13),.res(r27_14),.clk(clk),.wout(w27_14));
	PE pe27_15(.x(x15),.w(w27_14),.acc(r27_14),.res(r27_15),.clk(clk),.wout(w27_15));
	PE pe27_16(.x(x16),.w(w27_15),.acc(r27_15),.res(r27_16),.clk(clk),.wout(w27_16));
	PE pe27_17(.x(x17),.w(w27_16),.acc(r27_16),.res(r27_17),.clk(clk),.wout(w27_17));
	PE pe27_18(.x(x18),.w(w27_17),.acc(r27_17),.res(r27_18),.clk(clk),.wout(w27_18));
	PE pe27_19(.x(x19),.w(w27_18),.acc(r27_18),.res(r27_19),.clk(clk),.wout(w27_19));
	PE pe27_20(.x(x20),.w(w27_19),.acc(r27_19),.res(r27_20),.clk(clk),.wout(w27_20));
	PE pe27_21(.x(x21),.w(w27_20),.acc(r27_20),.res(r27_21),.clk(clk),.wout(w27_21));
	PE pe27_22(.x(x22),.w(w27_21),.acc(r27_21),.res(r27_22),.clk(clk),.wout(w27_22));
	PE pe27_23(.x(x23),.w(w27_22),.acc(r27_22),.res(r27_23),.clk(clk),.wout(w27_23));
	PE pe27_24(.x(x24),.w(w27_23),.acc(r27_23),.res(r27_24),.clk(clk),.wout(w27_24));
	PE pe27_25(.x(x25),.w(w27_24),.acc(r27_24),.res(r27_25),.clk(clk),.wout(w27_25));
	PE pe27_26(.x(x26),.w(w27_25),.acc(r27_25),.res(r27_26),.clk(clk),.wout(w27_26));
	PE pe27_27(.x(x27),.w(w27_26),.acc(r27_26),.res(r27_27),.clk(clk),.wout(w27_27));
	PE pe27_28(.x(x28),.w(w27_27),.acc(r27_27),.res(r27_28),.clk(clk),.wout(w27_28));
	PE pe27_29(.x(x29),.w(w27_28),.acc(r27_28),.res(r27_29),.clk(clk),.wout(w27_29));
	PE pe27_30(.x(x30),.w(w27_29),.acc(r27_29),.res(r27_30),.clk(clk),.wout(w27_30));
	PE pe27_31(.x(x31),.w(w27_30),.acc(r27_30),.res(r27_31),.clk(clk),.wout(w27_31));
	PE pe27_32(.x(x32),.w(w27_31),.acc(r27_31),.res(r27_32),.clk(clk),.wout(w27_32));
	PE pe27_33(.x(x33),.w(w27_32),.acc(r27_32),.res(r27_33),.clk(clk),.wout(w27_33));
	PE pe27_34(.x(x34),.w(w27_33),.acc(r27_33),.res(r27_34),.clk(clk),.wout(w27_34));
	PE pe27_35(.x(x35),.w(w27_34),.acc(r27_34),.res(r27_35),.clk(clk),.wout(w27_35));
	PE pe27_36(.x(x36),.w(w27_35),.acc(r27_35),.res(r27_36),.clk(clk),.wout(w27_36));
	PE pe27_37(.x(x37),.w(w27_36),.acc(r27_36),.res(r27_37),.clk(clk),.wout(w27_37));
	PE pe27_38(.x(x38),.w(w27_37),.acc(r27_37),.res(r27_38),.clk(clk),.wout(w27_38));
	PE pe27_39(.x(x39),.w(w27_38),.acc(r27_38),.res(r27_39),.clk(clk),.wout(w27_39));
	PE pe27_40(.x(x40),.w(w27_39),.acc(r27_39),.res(r27_40),.clk(clk),.wout(w27_40));
	PE pe27_41(.x(x41),.w(w27_40),.acc(r27_40),.res(r27_41),.clk(clk),.wout(w27_41));
	PE pe27_42(.x(x42),.w(w27_41),.acc(r27_41),.res(r27_42),.clk(clk),.wout(w27_42));
	PE pe27_43(.x(x43),.w(w27_42),.acc(r27_42),.res(r27_43),.clk(clk),.wout(w27_43));
	PE pe27_44(.x(x44),.w(w27_43),.acc(r27_43),.res(r27_44),.clk(clk),.wout(w27_44));
	PE pe27_45(.x(x45),.w(w27_44),.acc(r27_44),.res(r27_45),.clk(clk),.wout(w27_45));
	PE pe27_46(.x(x46),.w(w27_45),.acc(r27_45),.res(r27_46),.clk(clk),.wout(w27_46));
	PE pe27_47(.x(x47),.w(w27_46),.acc(r27_46),.res(r27_47),.clk(clk),.wout(w27_47));
	PE pe27_48(.x(x48),.w(w27_47),.acc(r27_47),.res(r27_48),.clk(clk),.wout(w27_48));
	PE pe27_49(.x(x49),.w(w27_48),.acc(r27_48),.res(r27_49),.clk(clk),.wout(w27_49));
	PE pe27_50(.x(x50),.w(w27_49),.acc(r27_49),.res(r27_50),.clk(clk),.wout(w27_50));
	PE pe27_51(.x(x51),.w(w27_50),.acc(r27_50),.res(r27_51),.clk(clk),.wout(w27_51));
	PE pe27_52(.x(x52),.w(w27_51),.acc(r27_51),.res(r27_52),.clk(clk),.wout(w27_52));
	PE pe27_53(.x(x53),.w(w27_52),.acc(r27_52),.res(r27_53),.clk(clk),.wout(w27_53));
	PE pe27_54(.x(x54),.w(w27_53),.acc(r27_53),.res(r27_54),.clk(clk),.wout(w27_54));
	PE pe27_55(.x(x55),.w(w27_54),.acc(r27_54),.res(r27_55),.clk(clk),.wout(w27_55));
	PE pe27_56(.x(x56),.w(w27_55),.acc(r27_55),.res(r27_56),.clk(clk),.wout(w27_56));
	PE pe27_57(.x(x57),.w(w27_56),.acc(r27_56),.res(r27_57),.clk(clk),.wout(w27_57));
	PE pe27_58(.x(x58),.w(w27_57),.acc(r27_57),.res(r27_58),.clk(clk),.wout(w27_58));
	PE pe27_59(.x(x59),.w(w27_58),.acc(r27_58),.res(r27_59),.clk(clk),.wout(w27_59));
	PE pe27_60(.x(x60),.w(w27_59),.acc(r27_59),.res(r27_60),.clk(clk),.wout(w27_60));
	PE pe27_61(.x(x61),.w(w27_60),.acc(r27_60),.res(r27_61),.clk(clk),.wout(w27_61));
	PE pe27_62(.x(x62),.w(w27_61),.acc(r27_61),.res(r27_62),.clk(clk),.wout(w27_62));
	PE pe27_63(.x(x63),.w(w27_62),.acc(r27_62),.res(r27_63),.clk(clk),.wout(w27_63));
	PE pe27_64(.x(x64),.w(w27_63),.acc(r27_63),.res(r27_64),.clk(clk),.wout(w27_64));
	PE pe27_65(.x(x65),.w(w27_64),.acc(r27_64),.res(r27_65),.clk(clk),.wout(w27_65));
	PE pe27_66(.x(x66),.w(w27_65),.acc(r27_65),.res(r27_66),.clk(clk),.wout(w27_66));
	PE pe27_67(.x(x67),.w(w27_66),.acc(r27_66),.res(r27_67),.clk(clk),.wout(w27_67));
	PE pe27_68(.x(x68),.w(w27_67),.acc(r27_67),.res(r27_68),.clk(clk),.wout(w27_68));
	PE pe27_69(.x(x69),.w(w27_68),.acc(r27_68),.res(r27_69),.clk(clk),.wout(w27_69));
	PE pe27_70(.x(x70),.w(w27_69),.acc(r27_69),.res(r27_70),.clk(clk),.wout(w27_70));
	PE pe27_71(.x(x71),.w(w27_70),.acc(r27_70),.res(r27_71),.clk(clk),.wout(w27_71));
	PE pe27_72(.x(x72),.w(w27_71),.acc(r27_71),.res(r27_72),.clk(clk),.wout(w27_72));
	PE pe27_73(.x(x73),.w(w27_72),.acc(r27_72),.res(r27_73),.clk(clk),.wout(w27_73));
	PE pe27_74(.x(x74),.w(w27_73),.acc(r27_73),.res(r27_74),.clk(clk),.wout(w27_74));
	PE pe27_75(.x(x75),.w(w27_74),.acc(r27_74),.res(r27_75),.clk(clk),.wout(w27_75));
	PE pe27_76(.x(x76),.w(w27_75),.acc(r27_75),.res(r27_76),.clk(clk),.wout(w27_76));
	PE pe27_77(.x(x77),.w(w27_76),.acc(r27_76),.res(r27_77),.clk(clk),.wout(w27_77));
	PE pe27_78(.x(x78),.w(w27_77),.acc(r27_77),.res(r27_78),.clk(clk),.wout(w27_78));
	PE pe27_79(.x(x79),.w(w27_78),.acc(r27_78),.res(r27_79),.clk(clk),.wout(w27_79));
	PE pe27_80(.x(x80),.w(w27_79),.acc(r27_79),.res(r27_80),.clk(clk),.wout(w27_80));
	PE pe27_81(.x(x81),.w(w27_80),.acc(r27_80),.res(r27_81),.clk(clk),.wout(w27_81));
	PE pe27_82(.x(x82),.w(w27_81),.acc(r27_81),.res(r27_82),.clk(clk),.wout(w27_82));
	PE pe27_83(.x(x83),.w(w27_82),.acc(r27_82),.res(r27_83),.clk(clk),.wout(w27_83));
	PE pe27_84(.x(x84),.w(w27_83),.acc(r27_83),.res(r27_84),.clk(clk),.wout(w27_84));
	PE pe27_85(.x(x85),.w(w27_84),.acc(r27_84),.res(r27_85),.clk(clk),.wout(w27_85));
	PE pe27_86(.x(x86),.w(w27_85),.acc(r27_85),.res(r27_86),.clk(clk),.wout(w27_86));
	PE pe27_87(.x(x87),.w(w27_86),.acc(r27_86),.res(r27_87),.clk(clk),.wout(w27_87));
	PE pe27_88(.x(x88),.w(w27_87),.acc(r27_87),.res(r27_88),.clk(clk),.wout(w27_88));
	PE pe27_89(.x(x89),.w(w27_88),.acc(r27_88),.res(r27_89),.clk(clk),.wout(w27_89));
	PE pe27_90(.x(x90),.w(w27_89),.acc(r27_89),.res(r27_90),.clk(clk),.wout(w27_90));
	PE pe27_91(.x(x91),.w(w27_90),.acc(r27_90),.res(r27_91),.clk(clk),.wout(w27_91));
	PE pe27_92(.x(x92),.w(w27_91),.acc(r27_91),.res(r27_92),.clk(clk),.wout(w27_92));
	PE pe27_93(.x(x93),.w(w27_92),.acc(r27_92),.res(r27_93),.clk(clk),.wout(w27_93));
	PE pe27_94(.x(x94),.w(w27_93),.acc(r27_93),.res(r27_94),.clk(clk),.wout(w27_94));
	PE pe27_95(.x(x95),.w(w27_94),.acc(r27_94),.res(r27_95),.clk(clk),.wout(w27_95));
	PE pe27_96(.x(x96),.w(w27_95),.acc(r27_95),.res(r27_96),.clk(clk),.wout(w27_96));
	PE pe27_97(.x(x97),.w(w27_96),.acc(r27_96),.res(r27_97),.clk(clk),.wout(w27_97));
	PE pe27_98(.x(x98),.w(w27_97),.acc(r27_97),.res(r27_98),.clk(clk),.wout(w27_98));
	PE pe27_99(.x(x99),.w(w27_98),.acc(r27_98),.res(r27_99),.clk(clk),.wout(w27_99));
	PE pe27_100(.x(x100),.w(w27_99),.acc(r27_99),.res(r27_100),.clk(clk),.wout(w27_100));
	PE pe27_101(.x(x101),.w(w27_100),.acc(r27_100),.res(r27_101),.clk(clk),.wout(w27_101));
	PE pe27_102(.x(x102),.w(w27_101),.acc(r27_101),.res(r27_102),.clk(clk),.wout(w27_102));
	PE pe27_103(.x(x103),.w(w27_102),.acc(r27_102),.res(r27_103),.clk(clk),.wout(w27_103));
	PE pe27_104(.x(x104),.w(w27_103),.acc(r27_103),.res(r27_104),.clk(clk),.wout(w27_104));
	PE pe27_105(.x(x105),.w(w27_104),.acc(r27_104),.res(r27_105),.clk(clk),.wout(w27_105));
	PE pe27_106(.x(x106),.w(w27_105),.acc(r27_105),.res(r27_106),.clk(clk),.wout(w27_106));
	PE pe27_107(.x(x107),.w(w27_106),.acc(r27_106),.res(r27_107),.clk(clk),.wout(w27_107));
	PE pe27_108(.x(x108),.w(w27_107),.acc(r27_107),.res(r27_108),.clk(clk),.wout(w27_108));
	PE pe27_109(.x(x109),.w(w27_108),.acc(r27_108),.res(r27_109),.clk(clk),.wout(w27_109));
	PE pe27_110(.x(x110),.w(w27_109),.acc(r27_109),.res(r27_110),.clk(clk),.wout(w27_110));
	PE pe27_111(.x(x111),.w(w27_110),.acc(r27_110),.res(r27_111),.clk(clk),.wout(w27_111));
	PE pe27_112(.x(x112),.w(w27_111),.acc(r27_111),.res(r27_112),.clk(clk),.wout(w27_112));
	PE pe27_113(.x(x113),.w(w27_112),.acc(r27_112),.res(r27_113),.clk(clk),.wout(w27_113));
	PE pe27_114(.x(x114),.w(w27_113),.acc(r27_113),.res(r27_114),.clk(clk),.wout(w27_114));
	PE pe27_115(.x(x115),.w(w27_114),.acc(r27_114),.res(r27_115),.clk(clk),.wout(w27_115));
	PE pe27_116(.x(x116),.w(w27_115),.acc(r27_115),.res(r27_116),.clk(clk),.wout(w27_116));
	PE pe27_117(.x(x117),.w(w27_116),.acc(r27_116),.res(r27_117),.clk(clk),.wout(w27_117));
	PE pe27_118(.x(x118),.w(w27_117),.acc(r27_117),.res(r27_118),.clk(clk),.wout(w27_118));
	PE pe27_119(.x(x119),.w(w27_118),.acc(r27_118),.res(r27_119),.clk(clk),.wout(w27_119));
	PE pe27_120(.x(x120),.w(w27_119),.acc(r27_119),.res(r27_120),.clk(clk),.wout(w27_120));
	PE pe27_121(.x(x121),.w(w27_120),.acc(r27_120),.res(r27_121),.clk(clk),.wout(w27_121));
	PE pe27_122(.x(x122),.w(w27_121),.acc(r27_121),.res(r27_122),.clk(clk),.wout(w27_122));
	PE pe27_123(.x(x123),.w(w27_122),.acc(r27_122),.res(r27_123),.clk(clk),.wout(w27_123));
	PE pe27_124(.x(x124),.w(w27_123),.acc(r27_123),.res(r27_124),.clk(clk),.wout(w27_124));
	PE pe27_125(.x(x125),.w(w27_124),.acc(r27_124),.res(r27_125),.clk(clk),.wout(w27_125));
	PE pe27_126(.x(x126),.w(w27_125),.acc(r27_125),.res(r27_126),.clk(clk),.wout(w27_126));
	PE pe27_127(.x(x127),.w(w27_126),.acc(r27_126),.res(result27),.clk(clk),.wout(weight27));

	PE pe28_0(.x(x0),.w(w28),.acc(32'h0),.res(r28_0),.clk(clk),.wout(w28_0));
	PE pe28_1(.x(x1),.w(w28_0),.acc(r28_0),.res(r28_1),.clk(clk),.wout(w28_1));
	PE pe28_2(.x(x2),.w(w28_1),.acc(r28_1),.res(r28_2),.clk(clk),.wout(w28_2));
	PE pe28_3(.x(x3),.w(w28_2),.acc(r28_2),.res(r28_3),.clk(clk),.wout(w28_3));
	PE pe28_4(.x(x4),.w(w28_3),.acc(r28_3),.res(r28_4),.clk(clk),.wout(w28_4));
	PE pe28_5(.x(x5),.w(w28_4),.acc(r28_4),.res(r28_5),.clk(clk),.wout(w28_5));
	PE pe28_6(.x(x6),.w(w28_5),.acc(r28_5),.res(r28_6),.clk(clk),.wout(w28_6));
	PE pe28_7(.x(x7),.w(w28_6),.acc(r28_6),.res(r28_7),.clk(clk),.wout(w28_7));
	PE pe28_8(.x(x8),.w(w28_7),.acc(r28_7),.res(r28_8),.clk(clk),.wout(w28_8));
	PE pe28_9(.x(x9),.w(w28_8),.acc(r28_8),.res(r28_9),.clk(clk),.wout(w28_9));
	PE pe28_10(.x(x10),.w(w28_9),.acc(r28_9),.res(r28_10),.clk(clk),.wout(w28_10));
	PE pe28_11(.x(x11),.w(w28_10),.acc(r28_10),.res(r28_11),.clk(clk),.wout(w28_11));
	PE pe28_12(.x(x12),.w(w28_11),.acc(r28_11),.res(r28_12),.clk(clk),.wout(w28_12));
	PE pe28_13(.x(x13),.w(w28_12),.acc(r28_12),.res(r28_13),.clk(clk),.wout(w28_13));
	PE pe28_14(.x(x14),.w(w28_13),.acc(r28_13),.res(r28_14),.clk(clk),.wout(w28_14));
	PE pe28_15(.x(x15),.w(w28_14),.acc(r28_14),.res(r28_15),.clk(clk),.wout(w28_15));
	PE pe28_16(.x(x16),.w(w28_15),.acc(r28_15),.res(r28_16),.clk(clk),.wout(w28_16));
	PE pe28_17(.x(x17),.w(w28_16),.acc(r28_16),.res(r28_17),.clk(clk),.wout(w28_17));
	PE pe28_18(.x(x18),.w(w28_17),.acc(r28_17),.res(r28_18),.clk(clk),.wout(w28_18));
	PE pe28_19(.x(x19),.w(w28_18),.acc(r28_18),.res(r28_19),.clk(clk),.wout(w28_19));
	PE pe28_20(.x(x20),.w(w28_19),.acc(r28_19),.res(r28_20),.clk(clk),.wout(w28_20));
	PE pe28_21(.x(x21),.w(w28_20),.acc(r28_20),.res(r28_21),.clk(clk),.wout(w28_21));
	PE pe28_22(.x(x22),.w(w28_21),.acc(r28_21),.res(r28_22),.clk(clk),.wout(w28_22));
	PE pe28_23(.x(x23),.w(w28_22),.acc(r28_22),.res(r28_23),.clk(clk),.wout(w28_23));
	PE pe28_24(.x(x24),.w(w28_23),.acc(r28_23),.res(r28_24),.clk(clk),.wout(w28_24));
	PE pe28_25(.x(x25),.w(w28_24),.acc(r28_24),.res(r28_25),.clk(clk),.wout(w28_25));
	PE pe28_26(.x(x26),.w(w28_25),.acc(r28_25),.res(r28_26),.clk(clk),.wout(w28_26));
	PE pe28_27(.x(x27),.w(w28_26),.acc(r28_26),.res(r28_27),.clk(clk),.wout(w28_27));
	PE pe28_28(.x(x28),.w(w28_27),.acc(r28_27),.res(r28_28),.clk(clk),.wout(w28_28));
	PE pe28_29(.x(x29),.w(w28_28),.acc(r28_28),.res(r28_29),.clk(clk),.wout(w28_29));
	PE pe28_30(.x(x30),.w(w28_29),.acc(r28_29),.res(r28_30),.clk(clk),.wout(w28_30));
	PE pe28_31(.x(x31),.w(w28_30),.acc(r28_30),.res(r28_31),.clk(clk),.wout(w28_31));
	PE pe28_32(.x(x32),.w(w28_31),.acc(r28_31),.res(r28_32),.clk(clk),.wout(w28_32));
	PE pe28_33(.x(x33),.w(w28_32),.acc(r28_32),.res(r28_33),.clk(clk),.wout(w28_33));
	PE pe28_34(.x(x34),.w(w28_33),.acc(r28_33),.res(r28_34),.clk(clk),.wout(w28_34));
	PE pe28_35(.x(x35),.w(w28_34),.acc(r28_34),.res(r28_35),.clk(clk),.wout(w28_35));
	PE pe28_36(.x(x36),.w(w28_35),.acc(r28_35),.res(r28_36),.clk(clk),.wout(w28_36));
	PE pe28_37(.x(x37),.w(w28_36),.acc(r28_36),.res(r28_37),.clk(clk),.wout(w28_37));
	PE pe28_38(.x(x38),.w(w28_37),.acc(r28_37),.res(r28_38),.clk(clk),.wout(w28_38));
	PE pe28_39(.x(x39),.w(w28_38),.acc(r28_38),.res(r28_39),.clk(clk),.wout(w28_39));
	PE pe28_40(.x(x40),.w(w28_39),.acc(r28_39),.res(r28_40),.clk(clk),.wout(w28_40));
	PE pe28_41(.x(x41),.w(w28_40),.acc(r28_40),.res(r28_41),.clk(clk),.wout(w28_41));
	PE pe28_42(.x(x42),.w(w28_41),.acc(r28_41),.res(r28_42),.clk(clk),.wout(w28_42));
	PE pe28_43(.x(x43),.w(w28_42),.acc(r28_42),.res(r28_43),.clk(clk),.wout(w28_43));
	PE pe28_44(.x(x44),.w(w28_43),.acc(r28_43),.res(r28_44),.clk(clk),.wout(w28_44));
	PE pe28_45(.x(x45),.w(w28_44),.acc(r28_44),.res(r28_45),.clk(clk),.wout(w28_45));
	PE pe28_46(.x(x46),.w(w28_45),.acc(r28_45),.res(r28_46),.clk(clk),.wout(w28_46));
	PE pe28_47(.x(x47),.w(w28_46),.acc(r28_46),.res(r28_47),.clk(clk),.wout(w28_47));
	PE pe28_48(.x(x48),.w(w28_47),.acc(r28_47),.res(r28_48),.clk(clk),.wout(w28_48));
	PE pe28_49(.x(x49),.w(w28_48),.acc(r28_48),.res(r28_49),.clk(clk),.wout(w28_49));
	PE pe28_50(.x(x50),.w(w28_49),.acc(r28_49),.res(r28_50),.clk(clk),.wout(w28_50));
	PE pe28_51(.x(x51),.w(w28_50),.acc(r28_50),.res(r28_51),.clk(clk),.wout(w28_51));
	PE pe28_52(.x(x52),.w(w28_51),.acc(r28_51),.res(r28_52),.clk(clk),.wout(w28_52));
	PE pe28_53(.x(x53),.w(w28_52),.acc(r28_52),.res(r28_53),.clk(clk),.wout(w28_53));
	PE pe28_54(.x(x54),.w(w28_53),.acc(r28_53),.res(r28_54),.clk(clk),.wout(w28_54));
	PE pe28_55(.x(x55),.w(w28_54),.acc(r28_54),.res(r28_55),.clk(clk),.wout(w28_55));
	PE pe28_56(.x(x56),.w(w28_55),.acc(r28_55),.res(r28_56),.clk(clk),.wout(w28_56));
	PE pe28_57(.x(x57),.w(w28_56),.acc(r28_56),.res(r28_57),.clk(clk),.wout(w28_57));
	PE pe28_58(.x(x58),.w(w28_57),.acc(r28_57),.res(r28_58),.clk(clk),.wout(w28_58));
	PE pe28_59(.x(x59),.w(w28_58),.acc(r28_58),.res(r28_59),.clk(clk),.wout(w28_59));
	PE pe28_60(.x(x60),.w(w28_59),.acc(r28_59),.res(r28_60),.clk(clk),.wout(w28_60));
	PE pe28_61(.x(x61),.w(w28_60),.acc(r28_60),.res(r28_61),.clk(clk),.wout(w28_61));
	PE pe28_62(.x(x62),.w(w28_61),.acc(r28_61),.res(r28_62),.clk(clk),.wout(w28_62));
	PE pe28_63(.x(x63),.w(w28_62),.acc(r28_62),.res(r28_63),.clk(clk),.wout(w28_63));
	PE pe28_64(.x(x64),.w(w28_63),.acc(r28_63),.res(r28_64),.clk(clk),.wout(w28_64));
	PE pe28_65(.x(x65),.w(w28_64),.acc(r28_64),.res(r28_65),.clk(clk),.wout(w28_65));
	PE pe28_66(.x(x66),.w(w28_65),.acc(r28_65),.res(r28_66),.clk(clk),.wout(w28_66));
	PE pe28_67(.x(x67),.w(w28_66),.acc(r28_66),.res(r28_67),.clk(clk),.wout(w28_67));
	PE pe28_68(.x(x68),.w(w28_67),.acc(r28_67),.res(r28_68),.clk(clk),.wout(w28_68));
	PE pe28_69(.x(x69),.w(w28_68),.acc(r28_68),.res(r28_69),.clk(clk),.wout(w28_69));
	PE pe28_70(.x(x70),.w(w28_69),.acc(r28_69),.res(r28_70),.clk(clk),.wout(w28_70));
	PE pe28_71(.x(x71),.w(w28_70),.acc(r28_70),.res(r28_71),.clk(clk),.wout(w28_71));
	PE pe28_72(.x(x72),.w(w28_71),.acc(r28_71),.res(r28_72),.clk(clk),.wout(w28_72));
	PE pe28_73(.x(x73),.w(w28_72),.acc(r28_72),.res(r28_73),.clk(clk),.wout(w28_73));
	PE pe28_74(.x(x74),.w(w28_73),.acc(r28_73),.res(r28_74),.clk(clk),.wout(w28_74));
	PE pe28_75(.x(x75),.w(w28_74),.acc(r28_74),.res(r28_75),.clk(clk),.wout(w28_75));
	PE pe28_76(.x(x76),.w(w28_75),.acc(r28_75),.res(r28_76),.clk(clk),.wout(w28_76));
	PE pe28_77(.x(x77),.w(w28_76),.acc(r28_76),.res(r28_77),.clk(clk),.wout(w28_77));
	PE pe28_78(.x(x78),.w(w28_77),.acc(r28_77),.res(r28_78),.clk(clk),.wout(w28_78));
	PE pe28_79(.x(x79),.w(w28_78),.acc(r28_78),.res(r28_79),.clk(clk),.wout(w28_79));
	PE pe28_80(.x(x80),.w(w28_79),.acc(r28_79),.res(r28_80),.clk(clk),.wout(w28_80));
	PE pe28_81(.x(x81),.w(w28_80),.acc(r28_80),.res(r28_81),.clk(clk),.wout(w28_81));
	PE pe28_82(.x(x82),.w(w28_81),.acc(r28_81),.res(r28_82),.clk(clk),.wout(w28_82));
	PE pe28_83(.x(x83),.w(w28_82),.acc(r28_82),.res(r28_83),.clk(clk),.wout(w28_83));
	PE pe28_84(.x(x84),.w(w28_83),.acc(r28_83),.res(r28_84),.clk(clk),.wout(w28_84));
	PE pe28_85(.x(x85),.w(w28_84),.acc(r28_84),.res(r28_85),.clk(clk),.wout(w28_85));
	PE pe28_86(.x(x86),.w(w28_85),.acc(r28_85),.res(r28_86),.clk(clk),.wout(w28_86));
	PE pe28_87(.x(x87),.w(w28_86),.acc(r28_86),.res(r28_87),.clk(clk),.wout(w28_87));
	PE pe28_88(.x(x88),.w(w28_87),.acc(r28_87),.res(r28_88),.clk(clk),.wout(w28_88));
	PE pe28_89(.x(x89),.w(w28_88),.acc(r28_88),.res(r28_89),.clk(clk),.wout(w28_89));
	PE pe28_90(.x(x90),.w(w28_89),.acc(r28_89),.res(r28_90),.clk(clk),.wout(w28_90));
	PE pe28_91(.x(x91),.w(w28_90),.acc(r28_90),.res(r28_91),.clk(clk),.wout(w28_91));
	PE pe28_92(.x(x92),.w(w28_91),.acc(r28_91),.res(r28_92),.clk(clk),.wout(w28_92));
	PE pe28_93(.x(x93),.w(w28_92),.acc(r28_92),.res(r28_93),.clk(clk),.wout(w28_93));
	PE pe28_94(.x(x94),.w(w28_93),.acc(r28_93),.res(r28_94),.clk(clk),.wout(w28_94));
	PE pe28_95(.x(x95),.w(w28_94),.acc(r28_94),.res(r28_95),.clk(clk),.wout(w28_95));
	PE pe28_96(.x(x96),.w(w28_95),.acc(r28_95),.res(r28_96),.clk(clk),.wout(w28_96));
	PE pe28_97(.x(x97),.w(w28_96),.acc(r28_96),.res(r28_97),.clk(clk),.wout(w28_97));
	PE pe28_98(.x(x98),.w(w28_97),.acc(r28_97),.res(r28_98),.clk(clk),.wout(w28_98));
	PE pe28_99(.x(x99),.w(w28_98),.acc(r28_98),.res(r28_99),.clk(clk),.wout(w28_99));
	PE pe28_100(.x(x100),.w(w28_99),.acc(r28_99),.res(r28_100),.clk(clk),.wout(w28_100));
	PE pe28_101(.x(x101),.w(w28_100),.acc(r28_100),.res(r28_101),.clk(clk),.wout(w28_101));
	PE pe28_102(.x(x102),.w(w28_101),.acc(r28_101),.res(r28_102),.clk(clk),.wout(w28_102));
	PE pe28_103(.x(x103),.w(w28_102),.acc(r28_102),.res(r28_103),.clk(clk),.wout(w28_103));
	PE pe28_104(.x(x104),.w(w28_103),.acc(r28_103),.res(r28_104),.clk(clk),.wout(w28_104));
	PE pe28_105(.x(x105),.w(w28_104),.acc(r28_104),.res(r28_105),.clk(clk),.wout(w28_105));
	PE pe28_106(.x(x106),.w(w28_105),.acc(r28_105),.res(r28_106),.clk(clk),.wout(w28_106));
	PE pe28_107(.x(x107),.w(w28_106),.acc(r28_106),.res(r28_107),.clk(clk),.wout(w28_107));
	PE pe28_108(.x(x108),.w(w28_107),.acc(r28_107),.res(r28_108),.clk(clk),.wout(w28_108));
	PE pe28_109(.x(x109),.w(w28_108),.acc(r28_108),.res(r28_109),.clk(clk),.wout(w28_109));
	PE pe28_110(.x(x110),.w(w28_109),.acc(r28_109),.res(r28_110),.clk(clk),.wout(w28_110));
	PE pe28_111(.x(x111),.w(w28_110),.acc(r28_110),.res(r28_111),.clk(clk),.wout(w28_111));
	PE pe28_112(.x(x112),.w(w28_111),.acc(r28_111),.res(r28_112),.clk(clk),.wout(w28_112));
	PE pe28_113(.x(x113),.w(w28_112),.acc(r28_112),.res(r28_113),.clk(clk),.wout(w28_113));
	PE pe28_114(.x(x114),.w(w28_113),.acc(r28_113),.res(r28_114),.clk(clk),.wout(w28_114));
	PE pe28_115(.x(x115),.w(w28_114),.acc(r28_114),.res(r28_115),.clk(clk),.wout(w28_115));
	PE pe28_116(.x(x116),.w(w28_115),.acc(r28_115),.res(r28_116),.clk(clk),.wout(w28_116));
	PE pe28_117(.x(x117),.w(w28_116),.acc(r28_116),.res(r28_117),.clk(clk),.wout(w28_117));
	PE pe28_118(.x(x118),.w(w28_117),.acc(r28_117),.res(r28_118),.clk(clk),.wout(w28_118));
	PE pe28_119(.x(x119),.w(w28_118),.acc(r28_118),.res(r28_119),.clk(clk),.wout(w28_119));
	PE pe28_120(.x(x120),.w(w28_119),.acc(r28_119),.res(r28_120),.clk(clk),.wout(w28_120));
	PE pe28_121(.x(x121),.w(w28_120),.acc(r28_120),.res(r28_121),.clk(clk),.wout(w28_121));
	PE pe28_122(.x(x122),.w(w28_121),.acc(r28_121),.res(r28_122),.clk(clk),.wout(w28_122));
	PE pe28_123(.x(x123),.w(w28_122),.acc(r28_122),.res(r28_123),.clk(clk),.wout(w28_123));
	PE pe28_124(.x(x124),.w(w28_123),.acc(r28_123),.res(r28_124),.clk(clk),.wout(w28_124));
	PE pe28_125(.x(x125),.w(w28_124),.acc(r28_124),.res(r28_125),.clk(clk),.wout(w28_125));
	PE pe28_126(.x(x126),.w(w28_125),.acc(r28_125),.res(r28_126),.clk(clk),.wout(w28_126));
	PE pe28_127(.x(x127),.w(w28_126),.acc(r28_126),.res(result28),.clk(clk),.wout(weight28));

	PE pe29_0(.x(x0),.w(w29),.acc(32'h0),.res(r29_0),.clk(clk),.wout(w29_0));
	PE pe29_1(.x(x1),.w(w29_0),.acc(r29_0),.res(r29_1),.clk(clk),.wout(w29_1));
	PE pe29_2(.x(x2),.w(w29_1),.acc(r29_1),.res(r29_2),.clk(clk),.wout(w29_2));
	PE pe29_3(.x(x3),.w(w29_2),.acc(r29_2),.res(r29_3),.clk(clk),.wout(w29_3));
	PE pe29_4(.x(x4),.w(w29_3),.acc(r29_3),.res(r29_4),.clk(clk),.wout(w29_4));
	PE pe29_5(.x(x5),.w(w29_4),.acc(r29_4),.res(r29_5),.clk(clk),.wout(w29_5));
	PE pe29_6(.x(x6),.w(w29_5),.acc(r29_5),.res(r29_6),.clk(clk),.wout(w29_6));
	PE pe29_7(.x(x7),.w(w29_6),.acc(r29_6),.res(r29_7),.clk(clk),.wout(w29_7));
	PE pe29_8(.x(x8),.w(w29_7),.acc(r29_7),.res(r29_8),.clk(clk),.wout(w29_8));
	PE pe29_9(.x(x9),.w(w29_8),.acc(r29_8),.res(r29_9),.clk(clk),.wout(w29_9));
	PE pe29_10(.x(x10),.w(w29_9),.acc(r29_9),.res(r29_10),.clk(clk),.wout(w29_10));
	PE pe29_11(.x(x11),.w(w29_10),.acc(r29_10),.res(r29_11),.clk(clk),.wout(w29_11));
	PE pe29_12(.x(x12),.w(w29_11),.acc(r29_11),.res(r29_12),.clk(clk),.wout(w29_12));
	PE pe29_13(.x(x13),.w(w29_12),.acc(r29_12),.res(r29_13),.clk(clk),.wout(w29_13));
	PE pe29_14(.x(x14),.w(w29_13),.acc(r29_13),.res(r29_14),.clk(clk),.wout(w29_14));
	PE pe29_15(.x(x15),.w(w29_14),.acc(r29_14),.res(r29_15),.clk(clk),.wout(w29_15));
	PE pe29_16(.x(x16),.w(w29_15),.acc(r29_15),.res(r29_16),.clk(clk),.wout(w29_16));
	PE pe29_17(.x(x17),.w(w29_16),.acc(r29_16),.res(r29_17),.clk(clk),.wout(w29_17));
	PE pe29_18(.x(x18),.w(w29_17),.acc(r29_17),.res(r29_18),.clk(clk),.wout(w29_18));
	PE pe29_19(.x(x19),.w(w29_18),.acc(r29_18),.res(r29_19),.clk(clk),.wout(w29_19));
	PE pe29_20(.x(x20),.w(w29_19),.acc(r29_19),.res(r29_20),.clk(clk),.wout(w29_20));
	PE pe29_21(.x(x21),.w(w29_20),.acc(r29_20),.res(r29_21),.clk(clk),.wout(w29_21));
	PE pe29_22(.x(x22),.w(w29_21),.acc(r29_21),.res(r29_22),.clk(clk),.wout(w29_22));
	PE pe29_23(.x(x23),.w(w29_22),.acc(r29_22),.res(r29_23),.clk(clk),.wout(w29_23));
	PE pe29_24(.x(x24),.w(w29_23),.acc(r29_23),.res(r29_24),.clk(clk),.wout(w29_24));
	PE pe29_25(.x(x25),.w(w29_24),.acc(r29_24),.res(r29_25),.clk(clk),.wout(w29_25));
	PE pe29_26(.x(x26),.w(w29_25),.acc(r29_25),.res(r29_26),.clk(clk),.wout(w29_26));
	PE pe29_27(.x(x27),.w(w29_26),.acc(r29_26),.res(r29_27),.clk(clk),.wout(w29_27));
	PE pe29_28(.x(x28),.w(w29_27),.acc(r29_27),.res(r29_28),.clk(clk),.wout(w29_28));
	PE pe29_29(.x(x29),.w(w29_28),.acc(r29_28),.res(r29_29),.clk(clk),.wout(w29_29));
	PE pe29_30(.x(x30),.w(w29_29),.acc(r29_29),.res(r29_30),.clk(clk),.wout(w29_30));
	PE pe29_31(.x(x31),.w(w29_30),.acc(r29_30),.res(r29_31),.clk(clk),.wout(w29_31));
	PE pe29_32(.x(x32),.w(w29_31),.acc(r29_31),.res(r29_32),.clk(clk),.wout(w29_32));
	PE pe29_33(.x(x33),.w(w29_32),.acc(r29_32),.res(r29_33),.clk(clk),.wout(w29_33));
	PE pe29_34(.x(x34),.w(w29_33),.acc(r29_33),.res(r29_34),.clk(clk),.wout(w29_34));
	PE pe29_35(.x(x35),.w(w29_34),.acc(r29_34),.res(r29_35),.clk(clk),.wout(w29_35));
	PE pe29_36(.x(x36),.w(w29_35),.acc(r29_35),.res(r29_36),.clk(clk),.wout(w29_36));
	PE pe29_37(.x(x37),.w(w29_36),.acc(r29_36),.res(r29_37),.clk(clk),.wout(w29_37));
	PE pe29_38(.x(x38),.w(w29_37),.acc(r29_37),.res(r29_38),.clk(clk),.wout(w29_38));
	PE pe29_39(.x(x39),.w(w29_38),.acc(r29_38),.res(r29_39),.clk(clk),.wout(w29_39));
	PE pe29_40(.x(x40),.w(w29_39),.acc(r29_39),.res(r29_40),.clk(clk),.wout(w29_40));
	PE pe29_41(.x(x41),.w(w29_40),.acc(r29_40),.res(r29_41),.clk(clk),.wout(w29_41));
	PE pe29_42(.x(x42),.w(w29_41),.acc(r29_41),.res(r29_42),.clk(clk),.wout(w29_42));
	PE pe29_43(.x(x43),.w(w29_42),.acc(r29_42),.res(r29_43),.clk(clk),.wout(w29_43));
	PE pe29_44(.x(x44),.w(w29_43),.acc(r29_43),.res(r29_44),.clk(clk),.wout(w29_44));
	PE pe29_45(.x(x45),.w(w29_44),.acc(r29_44),.res(r29_45),.clk(clk),.wout(w29_45));
	PE pe29_46(.x(x46),.w(w29_45),.acc(r29_45),.res(r29_46),.clk(clk),.wout(w29_46));
	PE pe29_47(.x(x47),.w(w29_46),.acc(r29_46),.res(r29_47),.clk(clk),.wout(w29_47));
	PE pe29_48(.x(x48),.w(w29_47),.acc(r29_47),.res(r29_48),.clk(clk),.wout(w29_48));
	PE pe29_49(.x(x49),.w(w29_48),.acc(r29_48),.res(r29_49),.clk(clk),.wout(w29_49));
	PE pe29_50(.x(x50),.w(w29_49),.acc(r29_49),.res(r29_50),.clk(clk),.wout(w29_50));
	PE pe29_51(.x(x51),.w(w29_50),.acc(r29_50),.res(r29_51),.clk(clk),.wout(w29_51));
	PE pe29_52(.x(x52),.w(w29_51),.acc(r29_51),.res(r29_52),.clk(clk),.wout(w29_52));
	PE pe29_53(.x(x53),.w(w29_52),.acc(r29_52),.res(r29_53),.clk(clk),.wout(w29_53));
	PE pe29_54(.x(x54),.w(w29_53),.acc(r29_53),.res(r29_54),.clk(clk),.wout(w29_54));
	PE pe29_55(.x(x55),.w(w29_54),.acc(r29_54),.res(r29_55),.clk(clk),.wout(w29_55));
	PE pe29_56(.x(x56),.w(w29_55),.acc(r29_55),.res(r29_56),.clk(clk),.wout(w29_56));
	PE pe29_57(.x(x57),.w(w29_56),.acc(r29_56),.res(r29_57),.clk(clk),.wout(w29_57));
	PE pe29_58(.x(x58),.w(w29_57),.acc(r29_57),.res(r29_58),.clk(clk),.wout(w29_58));
	PE pe29_59(.x(x59),.w(w29_58),.acc(r29_58),.res(r29_59),.clk(clk),.wout(w29_59));
	PE pe29_60(.x(x60),.w(w29_59),.acc(r29_59),.res(r29_60),.clk(clk),.wout(w29_60));
	PE pe29_61(.x(x61),.w(w29_60),.acc(r29_60),.res(r29_61),.clk(clk),.wout(w29_61));
	PE pe29_62(.x(x62),.w(w29_61),.acc(r29_61),.res(r29_62),.clk(clk),.wout(w29_62));
	PE pe29_63(.x(x63),.w(w29_62),.acc(r29_62),.res(r29_63),.clk(clk),.wout(w29_63));
	PE pe29_64(.x(x64),.w(w29_63),.acc(r29_63),.res(r29_64),.clk(clk),.wout(w29_64));
	PE pe29_65(.x(x65),.w(w29_64),.acc(r29_64),.res(r29_65),.clk(clk),.wout(w29_65));
	PE pe29_66(.x(x66),.w(w29_65),.acc(r29_65),.res(r29_66),.clk(clk),.wout(w29_66));
	PE pe29_67(.x(x67),.w(w29_66),.acc(r29_66),.res(r29_67),.clk(clk),.wout(w29_67));
	PE pe29_68(.x(x68),.w(w29_67),.acc(r29_67),.res(r29_68),.clk(clk),.wout(w29_68));
	PE pe29_69(.x(x69),.w(w29_68),.acc(r29_68),.res(r29_69),.clk(clk),.wout(w29_69));
	PE pe29_70(.x(x70),.w(w29_69),.acc(r29_69),.res(r29_70),.clk(clk),.wout(w29_70));
	PE pe29_71(.x(x71),.w(w29_70),.acc(r29_70),.res(r29_71),.clk(clk),.wout(w29_71));
	PE pe29_72(.x(x72),.w(w29_71),.acc(r29_71),.res(r29_72),.clk(clk),.wout(w29_72));
	PE pe29_73(.x(x73),.w(w29_72),.acc(r29_72),.res(r29_73),.clk(clk),.wout(w29_73));
	PE pe29_74(.x(x74),.w(w29_73),.acc(r29_73),.res(r29_74),.clk(clk),.wout(w29_74));
	PE pe29_75(.x(x75),.w(w29_74),.acc(r29_74),.res(r29_75),.clk(clk),.wout(w29_75));
	PE pe29_76(.x(x76),.w(w29_75),.acc(r29_75),.res(r29_76),.clk(clk),.wout(w29_76));
	PE pe29_77(.x(x77),.w(w29_76),.acc(r29_76),.res(r29_77),.clk(clk),.wout(w29_77));
	PE pe29_78(.x(x78),.w(w29_77),.acc(r29_77),.res(r29_78),.clk(clk),.wout(w29_78));
	PE pe29_79(.x(x79),.w(w29_78),.acc(r29_78),.res(r29_79),.clk(clk),.wout(w29_79));
	PE pe29_80(.x(x80),.w(w29_79),.acc(r29_79),.res(r29_80),.clk(clk),.wout(w29_80));
	PE pe29_81(.x(x81),.w(w29_80),.acc(r29_80),.res(r29_81),.clk(clk),.wout(w29_81));
	PE pe29_82(.x(x82),.w(w29_81),.acc(r29_81),.res(r29_82),.clk(clk),.wout(w29_82));
	PE pe29_83(.x(x83),.w(w29_82),.acc(r29_82),.res(r29_83),.clk(clk),.wout(w29_83));
	PE pe29_84(.x(x84),.w(w29_83),.acc(r29_83),.res(r29_84),.clk(clk),.wout(w29_84));
	PE pe29_85(.x(x85),.w(w29_84),.acc(r29_84),.res(r29_85),.clk(clk),.wout(w29_85));
	PE pe29_86(.x(x86),.w(w29_85),.acc(r29_85),.res(r29_86),.clk(clk),.wout(w29_86));
	PE pe29_87(.x(x87),.w(w29_86),.acc(r29_86),.res(r29_87),.clk(clk),.wout(w29_87));
	PE pe29_88(.x(x88),.w(w29_87),.acc(r29_87),.res(r29_88),.clk(clk),.wout(w29_88));
	PE pe29_89(.x(x89),.w(w29_88),.acc(r29_88),.res(r29_89),.clk(clk),.wout(w29_89));
	PE pe29_90(.x(x90),.w(w29_89),.acc(r29_89),.res(r29_90),.clk(clk),.wout(w29_90));
	PE pe29_91(.x(x91),.w(w29_90),.acc(r29_90),.res(r29_91),.clk(clk),.wout(w29_91));
	PE pe29_92(.x(x92),.w(w29_91),.acc(r29_91),.res(r29_92),.clk(clk),.wout(w29_92));
	PE pe29_93(.x(x93),.w(w29_92),.acc(r29_92),.res(r29_93),.clk(clk),.wout(w29_93));
	PE pe29_94(.x(x94),.w(w29_93),.acc(r29_93),.res(r29_94),.clk(clk),.wout(w29_94));
	PE pe29_95(.x(x95),.w(w29_94),.acc(r29_94),.res(r29_95),.clk(clk),.wout(w29_95));
	PE pe29_96(.x(x96),.w(w29_95),.acc(r29_95),.res(r29_96),.clk(clk),.wout(w29_96));
	PE pe29_97(.x(x97),.w(w29_96),.acc(r29_96),.res(r29_97),.clk(clk),.wout(w29_97));
	PE pe29_98(.x(x98),.w(w29_97),.acc(r29_97),.res(r29_98),.clk(clk),.wout(w29_98));
	PE pe29_99(.x(x99),.w(w29_98),.acc(r29_98),.res(r29_99),.clk(clk),.wout(w29_99));
	PE pe29_100(.x(x100),.w(w29_99),.acc(r29_99),.res(r29_100),.clk(clk),.wout(w29_100));
	PE pe29_101(.x(x101),.w(w29_100),.acc(r29_100),.res(r29_101),.clk(clk),.wout(w29_101));
	PE pe29_102(.x(x102),.w(w29_101),.acc(r29_101),.res(r29_102),.clk(clk),.wout(w29_102));
	PE pe29_103(.x(x103),.w(w29_102),.acc(r29_102),.res(r29_103),.clk(clk),.wout(w29_103));
	PE pe29_104(.x(x104),.w(w29_103),.acc(r29_103),.res(r29_104),.clk(clk),.wout(w29_104));
	PE pe29_105(.x(x105),.w(w29_104),.acc(r29_104),.res(r29_105),.clk(clk),.wout(w29_105));
	PE pe29_106(.x(x106),.w(w29_105),.acc(r29_105),.res(r29_106),.clk(clk),.wout(w29_106));
	PE pe29_107(.x(x107),.w(w29_106),.acc(r29_106),.res(r29_107),.clk(clk),.wout(w29_107));
	PE pe29_108(.x(x108),.w(w29_107),.acc(r29_107),.res(r29_108),.clk(clk),.wout(w29_108));
	PE pe29_109(.x(x109),.w(w29_108),.acc(r29_108),.res(r29_109),.clk(clk),.wout(w29_109));
	PE pe29_110(.x(x110),.w(w29_109),.acc(r29_109),.res(r29_110),.clk(clk),.wout(w29_110));
	PE pe29_111(.x(x111),.w(w29_110),.acc(r29_110),.res(r29_111),.clk(clk),.wout(w29_111));
	PE pe29_112(.x(x112),.w(w29_111),.acc(r29_111),.res(r29_112),.clk(clk),.wout(w29_112));
	PE pe29_113(.x(x113),.w(w29_112),.acc(r29_112),.res(r29_113),.clk(clk),.wout(w29_113));
	PE pe29_114(.x(x114),.w(w29_113),.acc(r29_113),.res(r29_114),.clk(clk),.wout(w29_114));
	PE pe29_115(.x(x115),.w(w29_114),.acc(r29_114),.res(r29_115),.clk(clk),.wout(w29_115));
	PE pe29_116(.x(x116),.w(w29_115),.acc(r29_115),.res(r29_116),.clk(clk),.wout(w29_116));
	PE pe29_117(.x(x117),.w(w29_116),.acc(r29_116),.res(r29_117),.clk(clk),.wout(w29_117));
	PE pe29_118(.x(x118),.w(w29_117),.acc(r29_117),.res(r29_118),.clk(clk),.wout(w29_118));
	PE pe29_119(.x(x119),.w(w29_118),.acc(r29_118),.res(r29_119),.clk(clk),.wout(w29_119));
	PE pe29_120(.x(x120),.w(w29_119),.acc(r29_119),.res(r29_120),.clk(clk),.wout(w29_120));
	PE pe29_121(.x(x121),.w(w29_120),.acc(r29_120),.res(r29_121),.clk(clk),.wout(w29_121));
	PE pe29_122(.x(x122),.w(w29_121),.acc(r29_121),.res(r29_122),.clk(clk),.wout(w29_122));
	PE pe29_123(.x(x123),.w(w29_122),.acc(r29_122),.res(r29_123),.clk(clk),.wout(w29_123));
	PE pe29_124(.x(x124),.w(w29_123),.acc(r29_123),.res(r29_124),.clk(clk),.wout(w29_124));
	PE pe29_125(.x(x125),.w(w29_124),.acc(r29_124),.res(r29_125),.clk(clk),.wout(w29_125));
	PE pe29_126(.x(x126),.w(w29_125),.acc(r29_125),.res(r29_126),.clk(clk),.wout(w29_126));
	PE pe29_127(.x(x127),.w(w29_126),.acc(r29_126),.res(result29),.clk(clk),.wout(weight29));

	PE pe30_0(.x(x0),.w(w30),.acc(32'h0),.res(r30_0),.clk(clk),.wout(w30_0));
	PE pe30_1(.x(x1),.w(w30_0),.acc(r30_0),.res(r30_1),.clk(clk),.wout(w30_1));
	PE pe30_2(.x(x2),.w(w30_1),.acc(r30_1),.res(r30_2),.clk(clk),.wout(w30_2));
	PE pe30_3(.x(x3),.w(w30_2),.acc(r30_2),.res(r30_3),.clk(clk),.wout(w30_3));
	PE pe30_4(.x(x4),.w(w30_3),.acc(r30_3),.res(r30_4),.clk(clk),.wout(w30_4));
	PE pe30_5(.x(x5),.w(w30_4),.acc(r30_4),.res(r30_5),.clk(clk),.wout(w30_5));
	PE pe30_6(.x(x6),.w(w30_5),.acc(r30_5),.res(r30_6),.clk(clk),.wout(w30_6));
	PE pe30_7(.x(x7),.w(w30_6),.acc(r30_6),.res(r30_7),.clk(clk),.wout(w30_7));
	PE pe30_8(.x(x8),.w(w30_7),.acc(r30_7),.res(r30_8),.clk(clk),.wout(w30_8));
	PE pe30_9(.x(x9),.w(w30_8),.acc(r30_8),.res(r30_9),.clk(clk),.wout(w30_9));
	PE pe30_10(.x(x10),.w(w30_9),.acc(r30_9),.res(r30_10),.clk(clk),.wout(w30_10));
	PE pe30_11(.x(x11),.w(w30_10),.acc(r30_10),.res(r30_11),.clk(clk),.wout(w30_11));
	PE pe30_12(.x(x12),.w(w30_11),.acc(r30_11),.res(r30_12),.clk(clk),.wout(w30_12));
	PE pe30_13(.x(x13),.w(w30_12),.acc(r30_12),.res(r30_13),.clk(clk),.wout(w30_13));
	PE pe30_14(.x(x14),.w(w30_13),.acc(r30_13),.res(r30_14),.clk(clk),.wout(w30_14));
	PE pe30_15(.x(x15),.w(w30_14),.acc(r30_14),.res(r30_15),.clk(clk),.wout(w30_15));
	PE pe30_16(.x(x16),.w(w30_15),.acc(r30_15),.res(r30_16),.clk(clk),.wout(w30_16));
	PE pe30_17(.x(x17),.w(w30_16),.acc(r30_16),.res(r30_17),.clk(clk),.wout(w30_17));
	PE pe30_18(.x(x18),.w(w30_17),.acc(r30_17),.res(r30_18),.clk(clk),.wout(w30_18));
	PE pe30_19(.x(x19),.w(w30_18),.acc(r30_18),.res(r30_19),.clk(clk),.wout(w30_19));
	PE pe30_20(.x(x20),.w(w30_19),.acc(r30_19),.res(r30_20),.clk(clk),.wout(w30_20));
	PE pe30_21(.x(x21),.w(w30_20),.acc(r30_20),.res(r30_21),.clk(clk),.wout(w30_21));
	PE pe30_22(.x(x22),.w(w30_21),.acc(r30_21),.res(r30_22),.clk(clk),.wout(w30_22));
	PE pe30_23(.x(x23),.w(w30_22),.acc(r30_22),.res(r30_23),.clk(clk),.wout(w30_23));
	PE pe30_24(.x(x24),.w(w30_23),.acc(r30_23),.res(r30_24),.clk(clk),.wout(w30_24));
	PE pe30_25(.x(x25),.w(w30_24),.acc(r30_24),.res(r30_25),.clk(clk),.wout(w30_25));
	PE pe30_26(.x(x26),.w(w30_25),.acc(r30_25),.res(r30_26),.clk(clk),.wout(w30_26));
	PE pe30_27(.x(x27),.w(w30_26),.acc(r30_26),.res(r30_27),.clk(clk),.wout(w30_27));
	PE pe30_28(.x(x28),.w(w30_27),.acc(r30_27),.res(r30_28),.clk(clk),.wout(w30_28));
	PE pe30_29(.x(x29),.w(w30_28),.acc(r30_28),.res(r30_29),.clk(clk),.wout(w30_29));
	PE pe30_30(.x(x30),.w(w30_29),.acc(r30_29),.res(r30_30),.clk(clk),.wout(w30_30));
	PE pe30_31(.x(x31),.w(w30_30),.acc(r30_30),.res(r30_31),.clk(clk),.wout(w30_31));
	PE pe30_32(.x(x32),.w(w30_31),.acc(r30_31),.res(r30_32),.clk(clk),.wout(w30_32));
	PE pe30_33(.x(x33),.w(w30_32),.acc(r30_32),.res(r30_33),.clk(clk),.wout(w30_33));
	PE pe30_34(.x(x34),.w(w30_33),.acc(r30_33),.res(r30_34),.clk(clk),.wout(w30_34));
	PE pe30_35(.x(x35),.w(w30_34),.acc(r30_34),.res(r30_35),.clk(clk),.wout(w30_35));
	PE pe30_36(.x(x36),.w(w30_35),.acc(r30_35),.res(r30_36),.clk(clk),.wout(w30_36));
	PE pe30_37(.x(x37),.w(w30_36),.acc(r30_36),.res(r30_37),.clk(clk),.wout(w30_37));
	PE pe30_38(.x(x38),.w(w30_37),.acc(r30_37),.res(r30_38),.clk(clk),.wout(w30_38));
	PE pe30_39(.x(x39),.w(w30_38),.acc(r30_38),.res(r30_39),.clk(clk),.wout(w30_39));
	PE pe30_40(.x(x40),.w(w30_39),.acc(r30_39),.res(r30_40),.clk(clk),.wout(w30_40));
	PE pe30_41(.x(x41),.w(w30_40),.acc(r30_40),.res(r30_41),.clk(clk),.wout(w30_41));
	PE pe30_42(.x(x42),.w(w30_41),.acc(r30_41),.res(r30_42),.clk(clk),.wout(w30_42));
	PE pe30_43(.x(x43),.w(w30_42),.acc(r30_42),.res(r30_43),.clk(clk),.wout(w30_43));
	PE pe30_44(.x(x44),.w(w30_43),.acc(r30_43),.res(r30_44),.clk(clk),.wout(w30_44));
	PE pe30_45(.x(x45),.w(w30_44),.acc(r30_44),.res(r30_45),.clk(clk),.wout(w30_45));
	PE pe30_46(.x(x46),.w(w30_45),.acc(r30_45),.res(r30_46),.clk(clk),.wout(w30_46));
	PE pe30_47(.x(x47),.w(w30_46),.acc(r30_46),.res(r30_47),.clk(clk),.wout(w30_47));
	PE pe30_48(.x(x48),.w(w30_47),.acc(r30_47),.res(r30_48),.clk(clk),.wout(w30_48));
	PE pe30_49(.x(x49),.w(w30_48),.acc(r30_48),.res(r30_49),.clk(clk),.wout(w30_49));
	PE pe30_50(.x(x50),.w(w30_49),.acc(r30_49),.res(r30_50),.clk(clk),.wout(w30_50));
	PE pe30_51(.x(x51),.w(w30_50),.acc(r30_50),.res(r30_51),.clk(clk),.wout(w30_51));
	PE pe30_52(.x(x52),.w(w30_51),.acc(r30_51),.res(r30_52),.clk(clk),.wout(w30_52));
	PE pe30_53(.x(x53),.w(w30_52),.acc(r30_52),.res(r30_53),.clk(clk),.wout(w30_53));
	PE pe30_54(.x(x54),.w(w30_53),.acc(r30_53),.res(r30_54),.clk(clk),.wout(w30_54));
	PE pe30_55(.x(x55),.w(w30_54),.acc(r30_54),.res(r30_55),.clk(clk),.wout(w30_55));
	PE pe30_56(.x(x56),.w(w30_55),.acc(r30_55),.res(r30_56),.clk(clk),.wout(w30_56));
	PE pe30_57(.x(x57),.w(w30_56),.acc(r30_56),.res(r30_57),.clk(clk),.wout(w30_57));
	PE pe30_58(.x(x58),.w(w30_57),.acc(r30_57),.res(r30_58),.clk(clk),.wout(w30_58));
	PE pe30_59(.x(x59),.w(w30_58),.acc(r30_58),.res(r30_59),.clk(clk),.wout(w30_59));
	PE pe30_60(.x(x60),.w(w30_59),.acc(r30_59),.res(r30_60),.clk(clk),.wout(w30_60));
	PE pe30_61(.x(x61),.w(w30_60),.acc(r30_60),.res(r30_61),.clk(clk),.wout(w30_61));
	PE pe30_62(.x(x62),.w(w30_61),.acc(r30_61),.res(r30_62),.clk(clk),.wout(w30_62));
	PE pe30_63(.x(x63),.w(w30_62),.acc(r30_62),.res(r30_63),.clk(clk),.wout(w30_63));
	PE pe30_64(.x(x64),.w(w30_63),.acc(r30_63),.res(r30_64),.clk(clk),.wout(w30_64));
	PE pe30_65(.x(x65),.w(w30_64),.acc(r30_64),.res(r30_65),.clk(clk),.wout(w30_65));
	PE pe30_66(.x(x66),.w(w30_65),.acc(r30_65),.res(r30_66),.clk(clk),.wout(w30_66));
	PE pe30_67(.x(x67),.w(w30_66),.acc(r30_66),.res(r30_67),.clk(clk),.wout(w30_67));
	PE pe30_68(.x(x68),.w(w30_67),.acc(r30_67),.res(r30_68),.clk(clk),.wout(w30_68));
	PE pe30_69(.x(x69),.w(w30_68),.acc(r30_68),.res(r30_69),.clk(clk),.wout(w30_69));
	PE pe30_70(.x(x70),.w(w30_69),.acc(r30_69),.res(r30_70),.clk(clk),.wout(w30_70));
	PE pe30_71(.x(x71),.w(w30_70),.acc(r30_70),.res(r30_71),.clk(clk),.wout(w30_71));
	PE pe30_72(.x(x72),.w(w30_71),.acc(r30_71),.res(r30_72),.clk(clk),.wout(w30_72));
	PE pe30_73(.x(x73),.w(w30_72),.acc(r30_72),.res(r30_73),.clk(clk),.wout(w30_73));
	PE pe30_74(.x(x74),.w(w30_73),.acc(r30_73),.res(r30_74),.clk(clk),.wout(w30_74));
	PE pe30_75(.x(x75),.w(w30_74),.acc(r30_74),.res(r30_75),.clk(clk),.wout(w30_75));
	PE pe30_76(.x(x76),.w(w30_75),.acc(r30_75),.res(r30_76),.clk(clk),.wout(w30_76));
	PE pe30_77(.x(x77),.w(w30_76),.acc(r30_76),.res(r30_77),.clk(clk),.wout(w30_77));
	PE pe30_78(.x(x78),.w(w30_77),.acc(r30_77),.res(r30_78),.clk(clk),.wout(w30_78));
	PE pe30_79(.x(x79),.w(w30_78),.acc(r30_78),.res(r30_79),.clk(clk),.wout(w30_79));
	PE pe30_80(.x(x80),.w(w30_79),.acc(r30_79),.res(r30_80),.clk(clk),.wout(w30_80));
	PE pe30_81(.x(x81),.w(w30_80),.acc(r30_80),.res(r30_81),.clk(clk),.wout(w30_81));
	PE pe30_82(.x(x82),.w(w30_81),.acc(r30_81),.res(r30_82),.clk(clk),.wout(w30_82));
	PE pe30_83(.x(x83),.w(w30_82),.acc(r30_82),.res(r30_83),.clk(clk),.wout(w30_83));
	PE pe30_84(.x(x84),.w(w30_83),.acc(r30_83),.res(r30_84),.clk(clk),.wout(w30_84));
	PE pe30_85(.x(x85),.w(w30_84),.acc(r30_84),.res(r30_85),.clk(clk),.wout(w30_85));
	PE pe30_86(.x(x86),.w(w30_85),.acc(r30_85),.res(r30_86),.clk(clk),.wout(w30_86));
	PE pe30_87(.x(x87),.w(w30_86),.acc(r30_86),.res(r30_87),.clk(clk),.wout(w30_87));
	PE pe30_88(.x(x88),.w(w30_87),.acc(r30_87),.res(r30_88),.clk(clk),.wout(w30_88));
	PE pe30_89(.x(x89),.w(w30_88),.acc(r30_88),.res(r30_89),.clk(clk),.wout(w30_89));
	PE pe30_90(.x(x90),.w(w30_89),.acc(r30_89),.res(r30_90),.clk(clk),.wout(w30_90));
	PE pe30_91(.x(x91),.w(w30_90),.acc(r30_90),.res(r30_91),.clk(clk),.wout(w30_91));
	PE pe30_92(.x(x92),.w(w30_91),.acc(r30_91),.res(r30_92),.clk(clk),.wout(w30_92));
	PE pe30_93(.x(x93),.w(w30_92),.acc(r30_92),.res(r30_93),.clk(clk),.wout(w30_93));
	PE pe30_94(.x(x94),.w(w30_93),.acc(r30_93),.res(r30_94),.clk(clk),.wout(w30_94));
	PE pe30_95(.x(x95),.w(w30_94),.acc(r30_94),.res(r30_95),.clk(clk),.wout(w30_95));
	PE pe30_96(.x(x96),.w(w30_95),.acc(r30_95),.res(r30_96),.clk(clk),.wout(w30_96));
	PE pe30_97(.x(x97),.w(w30_96),.acc(r30_96),.res(r30_97),.clk(clk),.wout(w30_97));
	PE pe30_98(.x(x98),.w(w30_97),.acc(r30_97),.res(r30_98),.clk(clk),.wout(w30_98));
	PE pe30_99(.x(x99),.w(w30_98),.acc(r30_98),.res(r30_99),.clk(clk),.wout(w30_99));
	PE pe30_100(.x(x100),.w(w30_99),.acc(r30_99),.res(r30_100),.clk(clk),.wout(w30_100));
	PE pe30_101(.x(x101),.w(w30_100),.acc(r30_100),.res(r30_101),.clk(clk),.wout(w30_101));
	PE pe30_102(.x(x102),.w(w30_101),.acc(r30_101),.res(r30_102),.clk(clk),.wout(w30_102));
	PE pe30_103(.x(x103),.w(w30_102),.acc(r30_102),.res(r30_103),.clk(clk),.wout(w30_103));
	PE pe30_104(.x(x104),.w(w30_103),.acc(r30_103),.res(r30_104),.clk(clk),.wout(w30_104));
	PE pe30_105(.x(x105),.w(w30_104),.acc(r30_104),.res(r30_105),.clk(clk),.wout(w30_105));
	PE pe30_106(.x(x106),.w(w30_105),.acc(r30_105),.res(r30_106),.clk(clk),.wout(w30_106));
	PE pe30_107(.x(x107),.w(w30_106),.acc(r30_106),.res(r30_107),.clk(clk),.wout(w30_107));
	PE pe30_108(.x(x108),.w(w30_107),.acc(r30_107),.res(r30_108),.clk(clk),.wout(w30_108));
	PE pe30_109(.x(x109),.w(w30_108),.acc(r30_108),.res(r30_109),.clk(clk),.wout(w30_109));
	PE pe30_110(.x(x110),.w(w30_109),.acc(r30_109),.res(r30_110),.clk(clk),.wout(w30_110));
	PE pe30_111(.x(x111),.w(w30_110),.acc(r30_110),.res(r30_111),.clk(clk),.wout(w30_111));
	PE pe30_112(.x(x112),.w(w30_111),.acc(r30_111),.res(r30_112),.clk(clk),.wout(w30_112));
	PE pe30_113(.x(x113),.w(w30_112),.acc(r30_112),.res(r30_113),.clk(clk),.wout(w30_113));
	PE pe30_114(.x(x114),.w(w30_113),.acc(r30_113),.res(r30_114),.clk(clk),.wout(w30_114));
	PE pe30_115(.x(x115),.w(w30_114),.acc(r30_114),.res(r30_115),.clk(clk),.wout(w30_115));
	PE pe30_116(.x(x116),.w(w30_115),.acc(r30_115),.res(r30_116),.clk(clk),.wout(w30_116));
	PE pe30_117(.x(x117),.w(w30_116),.acc(r30_116),.res(r30_117),.clk(clk),.wout(w30_117));
	PE pe30_118(.x(x118),.w(w30_117),.acc(r30_117),.res(r30_118),.clk(clk),.wout(w30_118));
	PE pe30_119(.x(x119),.w(w30_118),.acc(r30_118),.res(r30_119),.clk(clk),.wout(w30_119));
	PE pe30_120(.x(x120),.w(w30_119),.acc(r30_119),.res(r30_120),.clk(clk),.wout(w30_120));
	PE pe30_121(.x(x121),.w(w30_120),.acc(r30_120),.res(r30_121),.clk(clk),.wout(w30_121));
	PE pe30_122(.x(x122),.w(w30_121),.acc(r30_121),.res(r30_122),.clk(clk),.wout(w30_122));
	PE pe30_123(.x(x123),.w(w30_122),.acc(r30_122),.res(r30_123),.clk(clk),.wout(w30_123));
	PE pe30_124(.x(x124),.w(w30_123),.acc(r30_123),.res(r30_124),.clk(clk),.wout(w30_124));
	PE pe30_125(.x(x125),.w(w30_124),.acc(r30_124),.res(r30_125),.clk(clk),.wout(w30_125));
	PE pe30_126(.x(x126),.w(w30_125),.acc(r30_125),.res(r30_126),.clk(clk),.wout(w30_126));
	PE pe30_127(.x(x127),.w(w30_126),.acc(r30_126),.res(result30),.clk(clk),.wout(weight30));

	PE pe31_0(.x(x0),.w(w31),.acc(32'h0),.res(r31_0),.clk(clk),.wout(w31_0));
	PE pe31_1(.x(x1),.w(w31_0),.acc(r31_0),.res(r31_1),.clk(clk),.wout(w31_1));
	PE pe31_2(.x(x2),.w(w31_1),.acc(r31_1),.res(r31_2),.clk(clk),.wout(w31_2));
	PE pe31_3(.x(x3),.w(w31_2),.acc(r31_2),.res(r31_3),.clk(clk),.wout(w31_3));
	PE pe31_4(.x(x4),.w(w31_3),.acc(r31_3),.res(r31_4),.clk(clk),.wout(w31_4));
	PE pe31_5(.x(x5),.w(w31_4),.acc(r31_4),.res(r31_5),.clk(clk),.wout(w31_5));
	PE pe31_6(.x(x6),.w(w31_5),.acc(r31_5),.res(r31_6),.clk(clk),.wout(w31_6));
	PE pe31_7(.x(x7),.w(w31_6),.acc(r31_6),.res(r31_7),.clk(clk),.wout(w31_7));
	PE pe31_8(.x(x8),.w(w31_7),.acc(r31_7),.res(r31_8),.clk(clk),.wout(w31_8));
	PE pe31_9(.x(x9),.w(w31_8),.acc(r31_8),.res(r31_9),.clk(clk),.wout(w31_9));
	PE pe31_10(.x(x10),.w(w31_9),.acc(r31_9),.res(r31_10),.clk(clk),.wout(w31_10));
	PE pe31_11(.x(x11),.w(w31_10),.acc(r31_10),.res(r31_11),.clk(clk),.wout(w31_11));
	PE pe31_12(.x(x12),.w(w31_11),.acc(r31_11),.res(r31_12),.clk(clk),.wout(w31_12));
	PE pe31_13(.x(x13),.w(w31_12),.acc(r31_12),.res(r31_13),.clk(clk),.wout(w31_13));
	PE pe31_14(.x(x14),.w(w31_13),.acc(r31_13),.res(r31_14),.clk(clk),.wout(w31_14));
	PE pe31_15(.x(x15),.w(w31_14),.acc(r31_14),.res(r31_15),.clk(clk),.wout(w31_15));
	PE pe31_16(.x(x16),.w(w31_15),.acc(r31_15),.res(r31_16),.clk(clk),.wout(w31_16));
	PE pe31_17(.x(x17),.w(w31_16),.acc(r31_16),.res(r31_17),.clk(clk),.wout(w31_17));
	PE pe31_18(.x(x18),.w(w31_17),.acc(r31_17),.res(r31_18),.clk(clk),.wout(w31_18));
	PE pe31_19(.x(x19),.w(w31_18),.acc(r31_18),.res(r31_19),.clk(clk),.wout(w31_19));
	PE pe31_20(.x(x20),.w(w31_19),.acc(r31_19),.res(r31_20),.clk(clk),.wout(w31_20));
	PE pe31_21(.x(x21),.w(w31_20),.acc(r31_20),.res(r31_21),.clk(clk),.wout(w31_21));
	PE pe31_22(.x(x22),.w(w31_21),.acc(r31_21),.res(r31_22),.clk(clk),.wout(w31_22));
	PE pe31_23(.x(x23),.w(w31_22),.acc(r31_22),.res(r31_23),.clk(clk),.wout(w31_23));
	PE pe31_24(.x(x24),.w(w31_23),.acc(r31_23),.res(r31_24),.clk(clk),.wout(w31_24));
	PE pe31_25(.x(x25),.w(w31_24),.acc(r31_24),.res(r31_25),.clk(clk),.wout(w31_25));
	PE pe31_26(.x(x26),.w(w31_25),.acc(r31_25),.res(r31_26),.clk(clk),.wout(w31_26));
	PE pe31_27(.x(x27),.w(w31_26),.acc(r31_26),.res(r31_27),.clk(clk),.wout(w31_27));
	PE pe31_28(.x(x28),.w(w31_27),.acc(r31_27),.res(r31_28),.clk(clk),.wout(w31_28));
	PE pe31_29(.x(x29),.w(w31_28),.acc(r31_28),.res(r31_29),.clk(clk),.wout(w31_29));
	PE pe31_30(.x(x30),.w(w31_29),.acc(r31_29),.res(r31_30),.clk(clk),.wout(w31_30));
	PE pe31_31(.x(x31),.w(w31_30),.acc(r31_30),.res(r31_31),.clk(clk),.wout(w31_31));
	PE pe31_32(.x(x32),.w(w31_31),.acc(r31_31),.res(r31_32),.clk(clk),.wout(w31_32));
	PE pe31_33(.x(x33),.w(w31_32),.acc(r31_32),.res(r31_33),.clk(clk),.wout(w31_33));
	PE pe31_34(.x(x34),.w(w31_33),.acc(r31_33),.res(r31_34),.clk(clk),.wout(w31_34));
	PE pe31_35(.x(x35),.w(w31_34),.acc(r31_34),.res(r31_35),.clk(clk),.wout(w31_35));
	PE pe31_36(.x(x36),.w(w31_35),.acc(r31_35),.res(r31_36),.clk(clk),.wout(w31_36));
	PE pe31_37(.x(x37),.w(w31_36),.acc(r31_36),.res(r31_37),.clk(clk),.wout(w31_37));
	PE pe31_38(.x(x38),.w(w31_37),.acc(r31_37),.res(r31_38),.clk(clk),.wout(w31_38));
	PE pe31_39(.x(x39),.w(w31_38),.acc(r31_38),.res(r31_39),.clk(clk),.wout(w31_39));
	PE pe31_40(.x(x40),.w(w31_39),.acc(r31_39),.res(r31_40),.clk(clk),.wout(w31_40));
	PE pe31_41(.x(x41),.w(w31_40),.acc(r31_40),.res(r31_41),.clk(clk),.wout(w31_41));
	PE pe31_42(.x(x42),.w(w31_41),.acc(r31_41),.res(r31_42),.clk(clk),.wout(w31_42));
	PE pe31_43(.x(x43),.w(w31_42),.acc(r31_42),.res(r31_43),.clk(clk),.wout(w31_43));
	PE pe31_44(.x(x44),.w(w31_43),.acc(r31_43),.res(r31_44),.clk(clk),.wout(w31_44));
	PE pe31_45(.x(x45),.w(w31_44),.acc(r31_44),.res(r31_45),.clk(clk),.wout(w31_45));
	PE pe31_46(.x(x46),.w(w31_45),.acc(r31_45),.res(r31_46),.clk(clk),.wout(w31_46));
	PE pe31_47(.x(x47),.w(w31_46),.acc(r31_46),.res(r31_47),.clk(clk),.wout(w31_47));
	PE pe31_48(.x(x48),.w(w31_47),.acc(r31_47),.res(r31_48),.clk(clk),.wout(w31_48));
	PE pe31_49(.x(x49),.w(w31_48),.acc(r31_48),.res(r31_49),.clk(clk),.wout(w31_49));
	PE pe31_50(.x(x50),.w(w31_49),.acc(r31_49),.res(r31_50),.clk(clk),.wout(w31_50));
	PE pe31_51(.x(x51),.w(w31_50),.acc(r31_50),.res(r31_51),.clk(clk),.wout(w31_51));
	PE pe31_52(.x(x52),.w(w31_51),.acc(r31_51),.res(r31_52),.clk(clk),.wout(w31_52));
	PE pe31_53(.x(x53),.w(w31_52),.acc(r31_52),.res(r31_53),.clk(clk),.wout(w31_53));
	PE pe31_54(.x(x54),.w(w31_53),.acc(r31_53),.res(r31_54),.clk(clk),.wout(w31_54));
	PE pe31_55(.x(x55),.w(w31_54),.acc(r31_54),.res(r31_55),.clk(clk),.wout(w31_55));
	PE pe31_56(.x(x56),.w(w31_55),.acc(r31_55),.res(r31_56),.clk(clk),.wout(w31_56));
	PE pe31_57(.x(x57),.w(w31_56),.acc(r31_56),.res(r31_57),.clk(clk),.wout(w31_57));
	PE pe31_58(.x(x58),.w(w31_57),.acc(r31_57),.res(r31_58),.clk(clk),.wout(w31_58));
	PE pe31_59(.x(x59),.w(w31_58),.acc(r31_58),.res(r31_59),.clk(clk),.wout(w31_59));
	PE pe31_60(.x(x60),.w(w31_59),.acc(r31_59),.res(r31_60),.clk(clk),.wout(w31_60));
	PE pe31_61(.x(x61),.w(w31_60),.acc(r31_60),.res(r31_61),.clk(clk),.wout(w31_61));
	PE pe31_62(.x(x62),.w(w31_61),.acc(r31_61),.res(r31_62),.clk(clk),.wout(w31_62));
	PE pe31_63(.x(x63),.w(w31_62),.acc(r31_62),.res(r31_63),.clk(clk),.wout(w31_63));
	PE pe31_64(.x(x64),.w(w31_63),.acc(r31_63),.res(r31_64),.clk(clk),.wout(w31_64));
	PE pe31_65(.x(x65),.w(w31_64),.acc(r31_64),.res(r31_65),.clk(clk),.wout(w31_65));
	PE pe31_66(.x(x66),.w(w31_65),.acc(r31_65),.res(r31_66),.clk(clk),.wout(w31_66));
	PE pe31_67(.x(x67),.w(w31_66),.acc(r31_66),.res(r31_67),.clk(clk),.wout(w31_67));
	PE pe31_68(.x(x68),.w(w31_67),.acc(r31_67),.res(r31_68),.clk(clk),.wout(w31_68));
	PE pe31_69(.x(x69),.w(w31_68),.acc(r31_68),.res(r31_69),.clk(clk),.wout(w31_69));
	PE pe31_70(.x(x70),.w(w31_69),.acc(r31_69),.res(r31_70),.clk(clk),.wout(w31_70));
	PE pe31_71(.x(x71),.w(w31_70),.acc(r31_70),.res(r31_71),.clk(clk),.wout(w31_71));
	PE pe31_72(.x(x72),.w(w31_71),.acc(r31_71),.res(r31_72),.clk(clk),.wout(w31_72));
	PE pe31_73(.x(x73),.w(w31_72),.acc(r31_72),.res(r31_73),.clk(clk),.wout(w31_73));
	PE pe31_74(.x(x74),.w(w31_73),.acc(r31_73),.res(r31_74),.clk(clk),.wout(w31_74));
	PE pe31_75(.x(x75),.w(w31_74),.acc(r31_74),.res(r31_75),.clk(clk),.wout(w31_75));
	PE pe31_76(.x(x76),.w(w31_75),.acc(r31_75),.res(r31_76),.clk(clk),.wout(w31_76));
	PE pe31_77(.x(x77),.w(w31_76),.acc(r31_76),.res(r31_77),.clk(clk),.wout(w31_77));
	PE pe31_78(.x(x78),.w(w31_77),.acc(r31_77),.res(r31_78),.clk(clk),.wout(w31_78));
	PE pe31_79(.x(x79),.w(w31_78),.acc(r31_78),.res(r31_79),.clk(clk),.wout(w31_79));
	PE pe31_80(.x(x80),.w(w31_79),.acc(r31_79),.res(r31_80),.clk(clk),.wout(w31_80));
	PE pe31_81(.x(x81),.w(w31_80),.acc(r31_80),.res(r31_81),.clk(clk),.wout(w31_81));
	PE pe31_82(.x(x82),.w(w31_81),.acc(r31_81),.res(r31_82),.clk(clk),.wout(w31_82));
	PE pe31_83(.x(x83),.w(w31_82),.acc(r31_82),.res(r31_83),.clk(clk),.wout(w31_83));
	PE pe31_84(.x(x84),.w(w31_83),.acc(r31_83),.res(r31_84),.clk(clk),.wout(w31_84));
	PE pe31_85(.x(x85),.w(w31_84),.acc(r31_84),.res(r31_85),.clk(clk),.wout(w31_85));
	PE pe31_86(.x(x86),.w(w31_85),.acc(r31_85),.res(r31_86),.clk(clk),.wout(w31_86));
	PE pe31_87(.x(x87),.w(w31_86),.acc(r31_86),.res(r31_87),.clk(clk),.wout(w31_87));
	PE pe31_88(.x(x88),.w(w31_87),.acc(r31_87),.res(r31_88),.clk(clk),.wout(w31_88));
	PE pe31_89(.x(x89),.w(w31_88),.acc(r31_88),.res(r31_89),.clk(clk),.wout(w31_89));
	PE pe31_90(.x(x90),.w(w31_89),.acc(r31_89),.res(r31_90),.clk(clk),.wout(w31_90));
	PE pe31_91(.x(x91),.w(w31_90),.acc(r31_90),.res(r31_91),.clk(clk),.wout(w31_91));
	PE pe31_92(.x(x92),.w(w31_91),.acc(r31_91),.res(r31_92),.clk(clk),.wout(w31_92));
	PE pe31_93(.x(x93),.w(w31_92),.acc(r31_92),.res(r31_93),.clk(clk),.wout(w31_93));
	PE pe31_94(.x(x94),.w(w31_93),.acc(r31_93),.res(r31_94),.clk(clk),.wout(w31_94));
	PE pe31_95(.x(x95),.w(w31_94),.acc(r31_94),.res(r31_95),.clk(clk),.wout(w31_95));
	PE pe31_96(.x(x96),.w(w31_95),.acc(r31_95),.res(r31_96),.clk(clk),.wout(w31_96));
	PE pe31_97(.x(x97),.w(w31_96),.acc(r31_96),.res(r31_97),.clk(clk),.wout(w31_97));
	PE pe31_98(.x(x98),.w(w31_97),.acc(r31_97),.res(r31_98),.clk(clk),.wout(w31_98));
	PE pe31_99(.x(x99),.w(w31_98),.acc(r31_98),.res(r31_99),.clk(clk),.wout(w31_99));
	PE pe31_100(.x(x100),.w(w31_99),.acc(r31_99),.res(r31_100),.clk(clk),.wout(w31_100));
	PE pe31_101(.x(x101),.w(w31_100),.acc(r31_100),.res(r31_101),.clk(clk),.wout(w31_101));
	PE pe31_102(.x(x102),.w(w31_101),.acc(r31_101),.res(r31_102),.clk(clk),.wout(w31_102));
	PE pe31_103(.x(x103),.w(w31_102),.acc(r31_102),.res(r31_103),.clk(clk),.wout(w31_103));
	PE pe31_104(.x(x104),.w(w31_103),.acc(r31_103),.res(r31_104),.clk(clk),.wout(w31_104));
	PE pe31_105(.x(x105),.w(w31_104),.acc(r31_104),.res(r31_105),.clk(clk),.wout(w31_105));
	PE pe31_106(.x(x106),.w(w31_105),.acc(r31_105),.res(r31_106),.clk(clk),.wout(w31_106));
	PE pe31_107(.x(x107),.w(w31_106),.acc(r31_106),.res(r31_107),.clk(clk),.wout(w31_107));
	PE pe31_108(.x(x108),.w(w31_107),.acc(r31_107),.res(r31_108),.clk(clk),.wout(w31_108));
	PE pe31_109(.x(x109),.w(w31_108),.acc(r31_108),.res(r31_109),.clk(clk),.wout(w31_109));
	PE pe31_110(.x(x110),.w(w31_109),.acc(r31_109),.res(r31_110),.clk(clk),.wout(w31_110));
	PE pe31_111(.x(x111),.w(w31_110),.acc(r31_110),.res(r31_111),.clk(clk),.wout(w31_111));
	PE pe31_112(.x(x112),.w(w31_111),.acc(r31_111),.res(r31_112),.clk(clk),.wout(w31_112));
	PE pe31_113(.x(x113),.w(w31_112),.acc(r31_112),.res(r31_113),.clk(clk),.wout(w31_113));
	PE pe31_114(.x(x114),.w(w31_113),.acc(r31_113),.res(r31_114),.clk(clk),.wout(w31_114));
	PE pe31_115(.x(x115),.w(w31_114),.acc(r31_114),.res(r31_115),.clk(clk),.wout(w31_115));
	PE pe31_116(.x(x116),.w(w31_115),.acc(r31_115),.res(r31_116),.clk(clk),.wout(w31_116));
	PE pe31_117(.x(x117),.w(w31_116),.acc(r31_116),.res(r31_117),.clk(clk),.wout(w31_117));
	PE pe31_118(.x(x118),.w(w31_117),.acc(r31_117),.res(r31_118),.clk(clk),.wout(w31_118));
	PE pe31_119(.x(x119),.w(w31_118),.acc(r31_118),.res(r31_119),.clk(clk),.wout(w31_119));
	PE pe31_120(.x(x120),.w(w31_119),.acc(r31_119),.res(r31_120),.clk(clk),.wout(w31_120));
	PE pe31_121(.x(x121),.w(w31_120),.acc(r31_120),.res(r31_121),.clk(clk),.wout(w31_121));
	PE pe31_122(.x(x122),.w(w31_121),.acc(r31_121),.res(r31_122),.clk(clk),.wout(w31_122));
	PE pe31_123(.x(x123),.w(w31_122),.acc(r31_122),.res(r31_123),.clk(clk),.wout(w31_123));
	PE pe31_124(.x(x124),.w(w31_123),.acc(r31_123),.res(r31_124),.clk(clk),.wout(w31_124));
	PE pe31_125(.x(x125),.w(w31_124),.acc(r31_124),.res(r31_125),.clk(clk),.wout(w31_125));
	PE pe31_126(.x(x126),.w(w31_125),.acc(r31_125),.res(r31_126),.clk(clk),.wout(w31_126));
	PE pe31_127(.x(x127),.w(w31_126),.acc(r31_126),.res(result31),.clk(clk),.wout(weight31));

	PE pe32_0(.x(x0),.w(w32),.acc(32'h0),.res(r32_0),.clk(clk),.wout(w32_0));
	PE pe32_1(.x(x1),.w(w32_0),.acc(r32_0),.res(r32_1),.clk(clk),.wout(w32_1));
	PE pe32_2(.x(x2),.w(w32_1),.acc(r32_1),.res(r32_2),.clk(clk),.wout(w32_2));
	PE pe32_3(.x(x3),.w(w32_2),.acc(r32_2),.res(r32_3),.clk(clk),.wout(w32_3));
	PE pe32_4(.x(x4),.w(w32_3),.acc(r32_3),.res(r32_4),.clk(clk),.wout(w32_4));
	PE pe32_5(.x(x5),.w(w32_4),.acc(r32_4),.res(r32_5),.clk(clk),.wout(w32_5));
	PE pe32_6(.x(x6),.w(w32_5),.acc(r32_5),.res(r32_6),.clk(clk),.wout(w32_6));
	PE pe32_7(.x(x7),.w(w32_6),.acc(r32_6),.res(r32_7),.clk(clk),.wout(w32_7));
	PE pe32_8(.x(x8),.w(w32_7),.acc(r32_7),.res(r32_8),.clk(clk),.wout(w32_8));
	PE pe32_9(.x(x9),.w(w32_8),.acc(r32_8),.res(r32_9),.clk(clk),.wout(w32_9));
	PE pe32_10(.x(x10),.w(w32_9),.acc(r32_9),.res(r32_10),.clk(clk),.wout(w32_10));
	PE pe32_11(.x(x11),.w(w32_10),.acc(r32_10),.res(r32_11),.clk(clk),.wout(w32_11));
	PE pe32_12(.x(x12),.w(w32_11),.acc(r32_11),.res(r32_12),.clk(clk),.wout(w32_12));
	PE pe32_13(.x(x13),.w(w32_12),.acc(r32_12),.res(r32_13),.clk(clk),.wout(w32_13));
	PE pe32_14(.x(x14),.w(w32_13),.acc(r32_13),.res(r32_14),.clk(clk),.wout(w32_14));
	PE pe32_15(.x(x15),.w(w32_14),.acc(r32_14),.res(r32_15),.clk(clk),.wout(w32_15));
	PE pe32_16(.x(x16),.w(w32_15),.acc(r32_15),.res(r32_16),.clk(clk),.wout(w32_16));
	PE pe32_17(.x(x17),.w(w32_16),.acc(r32_16),.res(r32_17),.clk(clk),.wout(w32_17));
	PE pe32_18(.x(x18),.w(w32_17),.acc(r32_17),.res(r32_18),.clk(clk),.wout(w32_18));
	PE pe32_19(.x(x19),.w(w32_18),.acc(r32_18),.res(r32_19),.clk(clk),.wout(w32_19));
	PE pe32_20(.x(x20),.w(w32_19),.acc(r32_19),.res(r32_20),.clk(clk),.wout(w32_20));
	PE pe32_21(.x(x21),.w(w32_20),.acc(r32_20),.res(r32_21),.clk(clk),.wout(w32_21));
	PE pe32_22(.x(x22),.w(w32_21),.acc(r32_21),.res(r32_22),.clk(clk),.wout(w32_22));
	PE pe32_23(.x(x23),.w(w32_22),.acc(r32_22),.res(r32_23),.clk(clk),.wout(w32_23));
	PE pe32_24(.x(x24),.w(w32_23),.acc(r32_23),.res(r32_24),.clk(clk),.wout(w32_24));
	PE pe32_25(.x(x25),.w(w32_24),.acc(r32_24),.res(r32_25),.clk(clk),.wout(w32_25));
	PE pe32_26(.x(x26),.w(w32_25),.acc(r32_25),.res(r32_26),.clk(clk),.wout(w32_26));
	PE pe32_27(.x(x27),.w(w32_26),.acc(r32_26),.res(r32_27),.clk(clk),.wout(w32_27));
	PE pe32_28(.x(x28),.w(w32_27),.acc(r32_27),.res(r32_28),.clk(clk),.wout(w32_28));
	PE pe32_29(.x(x29),.w(w32_28),.acc(r32_28),.res(r32_29),.clk(clk),.wout(w32_29));
	PE pe32_30(.x(x30),.w(w32_29),.acc(r32_29),.res(r32_30),.clk(clk),.wout(w32_30));
	PE pe32_31(.x(x31),.w(w32_30),.acc(r32_30),.res(r32_31),.clk(clk),.wout(w32_31));
	PE pe32_32(.x(x32),.w(w32_31),.acc(r32_31),.res(r32_32),.clk(clk),.wout(w32_32));
	PE pe32_33(.x(x33),.w(w32_32),.acc(r32_32),.res(r32_33),.clk(clk),.wout(w32_33));
	PE pe32_34(.x(x34),.w(w32_33),.acc(r32_33),.res(r32_34),.clk(clk),.wout(w32_34));
	PE pe32_35(.x(x35),.w(w32_34),.acc(r32_34),.res(r32_35),.clk(clk),.wout(w32_35));
	PE pe32_36(.x(x36),.w(w32_35),.acc(r32_35),.res(r32_36),.clk(clk),.wout(w32_36));
	PE pe32_37(.x(x37),.w(w32_36),.acc(r32_36),.res(r32_37),.clk(clk),.wout(w32_37));
	PE pe32_38(.x(x38),.w(w32_37),.acc(r32_37),.res(r32_38),.clk(clk),.wout(w32_38));
	PE pe32_39(.x(x39),.w(w32_38),.acc(r32_38),.res(r32_39),.clk(clk),.wout(w32_39));
	PE pe32_40(.x(x40),.w(w32_39),.acc(r32_39),.res(r32_40),.clk(clk),.wout(w32_40));
	PE pe32_41(.x(x41),.w(w32_40),.acc(r32_40),.res(r32_41),.clk(clk),.wout(w32_41));
	PE pe32_42(.x(x42),.w(w32_41),.acc(r32_41),.res(r32_42),.clk(clk),.wout(w32_42));
	PE pe32_43(.x(x43),.w(w32_42),.acc(r32_42),.res(r32_43),.clk(clk),.wout(w32_43));
	PE pe32_44(.x(x44),.w(w32_43),.acc(r32_43),.res(r32_44),.clk(clk),.wout(w32_44));
	PE pe32_45(.x(x45),.w(w32_44),.acc(r32_44),.res(r32_45),.clk(clk),.wout(w32_45));
	PE pe32_46(.x(x46),.w(w32_45),.acc(r32_45),.res(r32_46),.clk(clk),.wout(w32_46));
	PE pe32_47(.x(x47),.w(w32_46),.acc(r32_46),.res(r32_47),.clk(clk),.wout(w32_47));
	PE pe32_48(.x(x48),.w(w32_47),.acc(r32_47),.res(r32_48),.clk(clk),.wout(w32_48));
	PE pe32_49(.x(x49),.w(w32_48),.acc(r32_48),.res(r32_49),.clk(clk),.wout(w32_49));
	PE pe32_50(.x(x50),.w(w32_49),.acc(r32_49),.res(r32_50),.clk(clk),.wout(w32_50));
	PE pe32_51(.x(x51),.w(w32_50),.acc(r32_50),.res(r32_51),.clk(clk),.wout(w32_51));
	PE pe32_52(.x(x52),.w(w32_51),.acc(r32_51),.res(r32_52),.clk(clk),.wout(w32_52));
	PE pe32_53(.x(x53),.w(w32_52),.acc(r32_52),.res(r32_53),.clk(clk),.wout(w32_53));
	PE pe32_54(.x(x54),.w(w32_53),.acc(r32_53),.res(r32_54),.clk(clk),.wout(w32_54));
	PE pe32_55(.x(x55),.w(w32_54),.acc(r32_54),.res(r32_55),.clk(clk),.wout(w32_55));
	PE pe32_56(.x(x56),.w(w32_55),.acc(r32_55),.res(r32_56),.clk(clk),.wout(w32_56));
	PE pe32_57(.x(x57),.w(w32_56),.acc(r32_56),.res(r32_57),.clk(clk),.wout(w32_57));
	PE pe32_58(.x(x58),.w(w32_57),.acc(r32_57),.res(r32_58),.clk(clk),.wout(w32_58));
	PE pe32_59(.x(x59),.w(w32_58),.acc(r32_58),.res(r32_59),.clk(clk),.wout(w32_59));
	PE pe32_60(.x(x60),.w(w32_59),.acc(r32_59),.res(r32_60),.clk(clk),.wout(w32_60));
	PE pe32_61(.x(x61),.w(w32_60),.acc(r32_60),.res(r32_61),.clk(clk),.wout(w32_61));
	PE pe32_62(.x(x62),.w(w32_61),.acc(r32_61),.res(r32_62),.clk(clk),.wout(w32_62));
	PE pe32_63(.x(x63),.w(w32_62),.acc(r32_62),.res(r32_63),.clk(clk),.wout(w32_63));
	PE pe32_64(.x(x64),.w(w32_63),.acc(r32_63),.res(r32_64),.clk(clk),.wout(w32_64));
	PE pe32_65(.x(x65),.w(w32_64),.acc(r32_64),.res(r32_65),.clk(clk),.wout(w32_65));
	PE pe32_66(.x(x66),.w(w32_65),.acc(r32_65),.res(r32_66),.clk(clk),.wout(w32_66));
	PE pe32_67(.x(x67),.w(w32_66),.acc(r32_66),.res(r32_67),.clk(clk),.wout(w32_67));
	PE pe32_68(.x(x68),.w(w32_67),.acc(r32_67),.res(r32_68),.clk(clk),.wout(w32_68));
	PE pe32_69(.x(x69),.w(w32_68),.acc(r32_68),.res(r32_69),.clk(clk),.wout(w32_69));
	PE pe32_70(.x(x70),.w(w32_69),.acc(r32_69),.res(r32_70),.clk(clk),.wout(w32_70));
	PE pe32_71(.x(x71),.w(w32_70),.acc(r32_70),.res(r32_71),.clk(clk),.wout(w32_71));
	PE pe32_72(.x(x72),.w(w32_71),.acc(r32_71),.res(r32_72),.clk(clk),.wout(w32_72));
	PE pe32_73(.x(x73),.w(w32_72),.acc(r32_72),.res(r32_73),.clk(clk),.wout(w32_73));
	PE pe32_74(.x(x74),.w(w32_73),.acc(r32_73),.res(r32_74),.clk(clk),.wout(w32_74));
	PE pe32_75(.x(x75),.w(w32_74),.acc(r32_74),.res(r32_75),.clk(clk),.wout(w32_75));
	PE pe32_76(.x(x76),.w(w32_75),.acc(r32_75),.res(r32_76),.clk(clk),.wout(w32_76));
	PE pe32_77(.x(x77),.w(w32_76),.acc(r32_76),.res(r32_77),.clk(clk),.wout(w32_77));
	PE pe32_78(.x(x78),.w(w32_77),.acc(r32_77),.res(r32_78),.clk(clk),.wout(w32_78));
	PE pe32_79(.x(x79),.w(w32_78),.acc(r32_78),.res(r32_79),.clk(clk),.wout(w32_79));
	PE pe32_80(.x(x80),.w(w32_79),.acc(r32_79),.res(r32_80),.clk(clk),.wout(w32_80));
	PE pe32_81(.x(x81),.w(w32_80),.acc(r32_80),.res(r32_81),.clk(clk),.wout(w32_81));
	PE pe32_82(.x(x82),.w(w32_81),.acc(r32_81),.res(r32_82),.clk(clk),.wout(w32_82));
	PE pe32_83(.x(x83),.w(w32_82),.acc(r32_82),.res(r32_83),.clk(clk),.wout(w32_83));
	PE pe32_84(.x(x84),.w(w32_83),.acc(r32_83),.res(r32_84),.clk(clk),.wout(w32_84));
	PE pe32_85(.x(x85),.w(w32_84),.acc(r32_84),.res(r32_85),.clk(clk),.wout(w32_85));
	PE pe32_86(.x(x86),.w(w32_85),.acc(r32_85),.res(r32_86),.clk(clk),.wout(w32_86));
	PE pe32_87(.x(x87),.w(w32_86),.acc(r32_86),.res(r32_87),.clk(clk),.wout(w32_87));
	PE pe32_88(.x(x88),.w(w32_87),.acc(r32_87),.res(r32_88),.clk(clk),.wout(w32_88));
	PE pe32_89(.x(x89),.w(w32_88),.acc(r32_88),.res(r32_89),.clk(clk),.wout(w32_89));
	PE pe32_90(.x(x90),.w(w32_89),.acc(r32_89),.res(r32_90),.clk(clk),.wout(w32_90));
	PE pe32_91(.x(x91),.w(w32_90),.acc(r32_90),.res(r32_91),.clk(clk),.wout(w32_91));
	PE pe32_92(.x(x92),.w(w32_91),.acc(r32_91),.res(r32_92),.clk(clk),.wout(w32_92));
	PE pe32_93(.x(x93),.w(w32_92),.acc(r32_92),.res(r32_93),.clk(clk),.wout(w32_93));
	PE pe32_94(.x(x94),.w(w32_93),.acc(r32_93),.res(r32_94),.clk(clk),.wout(w32_94));
	PE pe32_95(.x(x95),.w(w32_94),.acc(r32_94),.res(r32_95),.clk(clk),.wout(w32_95));
	PE pe32_96(.x(x96),.w(w32_95),.acc(r32_95),.res(r32_96),.clk(clk),.wout(w32_96));
	PE pe32_97(.x(x97),.w(w32_96),.acc(r32_96),.res(r32_97),.clk(clk),.wout(w32_97));
	PE pe32_98(.x(x98),.w(w32_97),.acc(r32_97),.res(r32_98),.clk(clk),.wout(w32_98));
	PE pe32_99(.x(x99),.w(w32_98),.acc(r32_98),.res(r32_99),.clk(clk),.wout(w32_99));
	PE pe32_100(.x(x100),.w(w32_99),.acc(r32_99),.res(r32_100),.clk(clk),.wout(w32_100));
	PE pe32_101(.x(x101),.w(w32_100),.acc(r32_100),.res(r32_101),.clk(clk),.wout(w32_101));
	PE pe32_102(.x(x102),.w(w32_101),.acc(r32_101),.res(r32_102),.clk(clk),.wout(w32_102));
	PE pe32_103(.x(x103),.w(w32_102),.acc(r32_102),.res(r32_103),.clk(clk),.wout(w32_103));
	PE pe32_104(.x(x104),.w(w32_103),.acc(r32_103),.res(r32_104),.clk(clk),.wout(w32_104));
	PE pe32_105(.x(x105),.w(w32_104),.acc(r32_104),.res(r32_105),.clk(clk),.wout(w32_105));
	PE pe32_106(.x(x106),.w(w32_105),.acc(r32_105),.res(r32_106),.clk(clk),.wout(w32_106));
	PE pe32_107(.x(x107),.w(w32_106),.acc(r32_106),.res(r32_107),.clk(clk),.wout(w32_107));
	PE pe32_108(.x(x108),.w(w32_107),.acc(r32_107),.res(r32_108),.clk(clk),.wout(w32_108));
	PE pe32_109(.x(x109),.w(w32_108),.acc(r32_108),.res(r32_109),.clk(clk),.wout(w32_109));
	PE pe32_110(.x(x110),.w(w32_109),.acc(r32_109),.res(r32_110),.clk(clk),.wout(w32_110));
	PE pe32_111(.x(x111),.w(w32_110),.acc(r32_110),.res(r32_111),.clk(clk),.wout(w32_111));
	PE pe32_112(.x(x112),.w(w32_111),.acc(r32_111),.res(r32_112),.clk(clk),.wout(w32_112));
	PE pe32_113(.x(x113),.w(w32_112),.acc(r32_112),.res(r32_113),.clk(clk),.wout(w32_113));
	PE pe32_114(.x(x114),.w(w32_113),.acc(r32_113),.res(r32_114),.clk(clk),.wout(w32_114));
	PE pe32_115(.x(x115),.w(w32_114),.acc(r32_114),.res(r32_115),.clk(clk),.wout(w32_115));
	PE pe32_116(.x(x116),.w(w32_115),.acc(r32_115),.res(r32_116),.clk(clk),.wout(w32_116));
	PE pe32_117(.x(x117),.w(w32_116),.acc(r32_116),.res(r32_117),.clk(clk),.wout(w32_117));
	PE pe32_118(.x(x118),.w(w32_117),.acc(r32_117),.res(r32_118),.clk(clk),.wout(w32_118));
	PE pe32_119(.x(x119),.w(w32_118),.acc(r32_118),.res(r32_119),.clk(clk),.wout(w32_119));
	PE pe32_120(.x(x120),.w(w32_119),.acc(r32_119),.res(r32_120),.clk(clk),.wout(w32_120));
	PE pe32_121(.x(x121),.w(w32_120),.acc(r32_120),.res(r32_121),.clk(clk),.wout(w32_121));
	PE pe32_122(.x(x122),.w(w32_121),.acc(r32_121),.res(r32_122),.clk(clk),.wout(w32_122));
	PE pe32_123(.x(x123),.w(w32_122),.acc(r32_122),.res(r32_123),.clk(clk),.wout(w32_123));
	PE pe32_124(.x(x124),.w(w32_123),.acc(r32_123),.res(r32_124),.clk(clk),.wout(w32_124));
	PE pe32_125(.x(x125),.w(w32_124),.acc(r32_124),.res(r32_125),.clk(clk),.wout(w32_125));
	PE pe32_126(.x(x126),.w(w32_125),.acc(r32_125),.res(r32_126),.clk(clk),.wout(w32_126));
	PE pe32_127(.x(x127),.w(w32_126),.acc(r32_126),.res(result32),.clk(clk),.wout(weight32));

	PE pe33_0(.x(x0),.w(w33),.acc(32'h0),.res(r33_0),.clk(clk),.wout(w33_0));
	PE pe33_1(.x(x1),.w(w33_0),.acc(r33_0),.res(r33_1),.clk(clk),.wout(w33_1));
	PE pe33_2(.x(x2),.w(w33_1),.acc(r33_1),.res(r33_2),.clk(clk),.wout(w33_2));
	PE pe33_3(.x(x3),.w(w33_2),.acc(r33_2),.res(r33_3),.clk(clk),.wout(w33_3));
	PE pe33_4(.x(x4),.w(w33_3),.acc(r33_3),.res(r33_4),.clk(clk),.wout(w33_4));
	PE pe33_5(.x(x5),.w(w33_4),.acc(r33_4),.res(r33_5),.clk(clk),.wout(w33_5));
	PE pe33_6(.x(x6),.w(w33_5),.acc(r33_5),.res(r33_6),.clk(clk),.wout(w33_6));
	PE pe33_7(.x(x7),.w(w33_6),.acc(r33_6),.res(r33_7),.clk(clk),.wout(w33_7));
	PE pe33_8(.x(x8),.w(w33_7),.acc(r33_7),.res(r33_8),.clk(clk),.wout(w33_8));
	PE pe33_9(.x(x9),.w(w33_8),.acc(r33_8),.res(r33_9),.clk(clk),.wout(w33_9));
	PE pe33_10(.x(x10),.w(w33_9),.acc(r33_9),.res(r33_10),.clk(clk),.wout(w33_10));
	PE pe33_11(.x(x11),.w(w33_10),.acc(r33_10),.res(r33_11),.clk(clk),.wout(w33_11));
	PE pe33_12(.x(x12),.w(w33_11),.acc(r33_11),.res(r33_12),.clk(clk),.wout(w33_12));
	PE pe33_13(.x(x13),.w(w33_12),.acc(r33_12),.res(r33_13),.clk(clk),.wout(w33_13));
	PE pe33_14(.x(x14),.w(w33_13),.acc(r33_13),.res(r33_14),.clk(clk),.wout(w33_14));
	PE pe33_15(.x(x15),.w(w33_14),.acc(r33_14),.res(r33_15),.clk(clk),.wout(w33_15));
	PE pe33_16(.x(x16),.w(w33_15),.acc(r33_15),.res(r33_16),.clk(clk),.wout(w33_16));
	PE pe33_17(.x(x17),.w(w33_16),.acc(r33_16),.res(r33_17),.clk(clk),.wout(w33_17));
	PE pe33_18(.x(x18),.w(w33_17),.acc(r33_17),.res(r33_18),.clk(clk),.wout(w33_18));
	PE pe33_19(.x(x19),.w(w33_18),.acc(r33_18),.res(r33_19),.clk(clk),.wout(w33_19));
	PE pe33_20(.x(x20),.w(w33_19),.acc(r33_19),.res(r33_20),.clk(clk),.wout(w33_20));
	PE pe33_21(.x(x21),.w(w33_20),.acc(r33_20),.res(r33_21),.clk(clk),.wout(w33_21));
	PE pe33_22(.x(x22),.w(w33_21),.acc(r33_21),.res(r33_22),.clk(clk),.wout(w33_22));
	PE pe33_23(.x(x23),.w(w33_22),.acc(r33_22),.res(r33_23),.clk(clk),.wout(w33_23));
	PE pe33_24(.x(x24),.w(w33_23),.acc(r33_23),.res(r33_24),.clk(clk),.wout(w33_24));
	PE pe33_25(.x(x25),.w(w33_24),.acc(r33_24),.res(r33_25),.clk(clk),.wout(w33_25));
	PE pe33_26(.x(x26),.w(w33_25),.acc(r33_25),.res(r33_26),.clk(clk),.wout(w33_26));
	PE pe33_27(.x(x27),.w(w33_26),.acc(r33_26),.res(r33_27),.clk(clk),.wout(w33_27));
	PE pe33_28(.x(x28),.w(w33_27),.acc(r33_27),.res(r33_28),.clk(clk),.wout(w33_28));
	PE pe33_29(.x(x29),.w(w33_28),.acc(r33_28),.res(r33_29),.clk(clk),.wout(w33_29));
	PE pe33_30(.x(x30),.w(w33_29),.acc(r33_29),.res(r33_30),.clk(clk),.wout(w33_30));
	PE pe33_31(.x(x31),.w(w33_30),.acc(r33_30),.res(r33_31),.clk(clk),.wout(w33_31));
	PE pe33_32(.x(x32),.w(w33_31),.acc(r33_31),.res(r33_32),.clk(clk),.wout(w33_32));
	PE pe33_33(.x(x33),.w(w33_32),.acc(r33_32),.res(r33_33),.clk(clk),.wout(w33_33));
	PE pe33_34(.x(x34),.w(w33_33),.acc(r33_33),.res(r33_34),.clk(clk),.wout(w33_34));
	PE pe33_35(.x(x35),.w(w33_34),.acc(r33_34),.res(r33_35),.clk(clk),.wout(w33_35));
	PE pe33_36(.x(x36),.w(w33_35),.acc(r33_35),.res(r33_36),.clk(clk),.wout(w33_36));
	PE pe33_37(.x(x37),.w(w33_36),.acc(r33_36),.res(r33_37),.clk(clk),.wout(w33_37));
	PE pe33_38(.x(x38),.w(w33_37),.acc(r33_37),.res(r33_38),.clk(clk),.wout(w33_38));
	PE pe33_39(.x(x39),.w(w33_38),.acc(r33_38),.res(r33_39),.clk(clk),.wout(w33_39));
	PE pe33_40(.x(x40),.w(w33_39),.acc(r33_39),.res(r33_40),.clk(clk),.wout(w33_40));
	PE pe33_41(.x(x41),.w(w33_40),.acc(r33_40),.res(r33_41),.clk(clk),.wout(w33_41));
	PE pe33_42(.x(x42),.w(w33_41),.acc(r33_41),.res(r33_42),.clk(clk),.wout(w33_42));
	PE pe33_43(.x(x43),.w(w33_42),.acc(r33_42),.res(r33_43),.clk(clk),.wout(w33_43));
	PE pe33_44(.x(x44),.w(w33_43),.acc(r33_43),.res(r33_44),.clk(clk),.wout(w33_44));
	PE pe33_45(.x(x45),.w(w33_44),.acc(r33_44),.res(r33_45),.clk(clk),.wout(w33_45));
	PE pe33_46(.x(x46),.w(w33_45),.acc(r33_45),.res(r33_46),.clk(clk),.wout(w33_46));
	PE pe33_47(.x(x47),.w(w33_46),.acc(r33_46),.res(r33_47),.clk(clk),.wout(w33_47));
	PE pe33_48(.x(x48),.w(w33_47),.acc(r33_47),.res(r33_48),.clk(clk),.wout(w33_48));
	PE pe33_49(.x(x49),.w(w33_48),.acc(r33_48),.res(r33_49),.clk(clk),.wout(w33_49));
	PE pe33_50(.x(x50),.w(w33_49),.acc(r33_49),.res(r33_50),.clk(clk),.wout(w33_50));
	PE pe33_51(.x(x51),.w(w33_50),.acc(r33_50),.res(r33_51),.clk(clk),.wout(w33_51));
	PE pe33_52(.x(x52),.w(w33_51),.acc(r33_51),.res(r33_52),.clk(clk),.wout(w33_52));
	PE pe33_53(.x(x53),.w(w33_52),.acc(r33_52),.res(r33_53),.clk(clk),.wout(w33_53));
	PE pe33_54(.x(x54),.w(w33_53),.acc(r33_53),.res(r33_54),.clk(clk),.wout(w33_54));
	PE pe33_55(.x(x55),.w(w33_54),.acc(r33_54),.res(r33_55),.clk(clk),.wout(w33_55));
	PE pe33_56(.x(x56),.w(w33_55),.acc(r33_55),.res(r33_56),.clk(clk),.wout(w33_56));
	PE pe33_57(.x(x57),.w(w33_56),.acc(r33_56),.res(r33_57),.clk(clk),.wout(w33_57));
	PE pe33_58(.x(x58),.w(w33_57),.acc(r33_57),.res(r33_58),.clk(clk),.wout(w33_58));
	PE pe33_59(.x(x59),.w(w33_58),.acc(r33_58),.res(r33_59),.clk(clk),.wout(w33_59));
	PE pe33_60(.x(x60),.w(w33_59),.acc(r33_59),.res(r33_60),.clk(clk),.wout(w33_60));
	PE pe33_61(.x(x61),.w(w33_60),.acc(r33_60),.res(r33_61),.clk(clk),.wout(w33_61));
	PE pe33_62(.x(x62),.w(w33_61),.acc(r33_61),.res(r33_62),.clk(clk),.wout(w33_62));
	PE pe33_63(.x(x63),.w(w33_62),.acc(r33_62),.res(r33_63),.clk(clk),.wout(w33_63));
	PE pe33_64(.x(x64),.w(w33_63),.acc(r33_63),.res(r33_64),.clk(clk),.wout(w33_64));
	PE pe33_65(.x(x65),.w(w33_64),.acc(r33_64),.res(r33_65),.clk(clk),.wout(w33_65));
	PE pe33_66(.x(x66),.w(w33_65),.acc(r33_65),.res(r33_66),.clk(clk),.wout(w33_66));
	PE pe33_67(.x(x67),.w(w33_66),.acc(r33_66),.res(r33_67),.clk(clk),.wout(w33_67));
	PE pe33_68(.x(x68),.w(w33_67),.acc(r33_67),.res(r33_68),.clk(clk),.wout(w33_68));
	PE pe33_69(.x(x69),.w(w33_68),.acc(r33_68),.res(r33_69),.clk(clk),.wout(w33_69));
	PE pe33_70(.x(x70),.w(w33_69),.acc(r33_69),.res(r33_70),.clk(clk),.wout(w33_70));
	PE pe33_71(.x(x71),.w(w33_70),.acc(r33_70),.res(r33_71),.clk(clk),.wout(w33_71));
	PE pe33_72(.x(x72),.w(w33_71),.acc(r33_71),.res(r33_72),.clk(clk),.wout(w33_72));
	PE pe33_73(.x(x73),.w(w33_72),.acc(r33_72),.res(r33_73),.clk(clk),.wout(w33_73));
	PE pe33_74(.x(x74),.w(w33_73),.acc(r33_73),.res(r33_74),.clk(clk),.wout(w33_74));
	PE pe33_75(.x(x75),.w(w33_74),.acc(r33_74),.res(r33_75),.clk(clk),.wout(w33_75));
	PE pe33_76(.x(x76),.w(w33_75),.acc(r33_75),.res(r33_76),.clk(clk),.wout(w33_76));
	PE pe33_77(.x(x77),.w(w33_76),.acc(r33_76),.res(r33_77),.clk(clk),.wout(w33_77));
	PE pe33_78(.x(x78),.w(w33_77),.acc(r33_77),.res(r33_78),.clk(clk),.wout(w33_78));
	PE pe33_79(.x(x79),.w(w33_78),.acc(r33_78),.res(r33_79),.clk(clk),.wout(w33_79));
	PE pe33_80(.x(x80),.w(w33_79),.acc(r33_79),.res(r33_80),.clk(clk),.wout(w33_80));
	PE pe33_81(.x(x81),.w(w33_80),.acc(r33_80),.res(r33_81),.clk(clk),.wout(w33_81));
	PE pe33_82(.x(x82),.w(w33_81),.acc(r33_81),.res(r33_82),.clk(clk),.wout(w33_82));
	PE pe33_83(.x(x83),.w(w33_82),.acc(r33_82),.res(r33_83),.clk(clk),.wout(w33_83));
	PE pe33_84(.x(x84),.w(w33_83),.acc(r33_83),.res(r33_84),.clk(clk),.wout(w33_84));
	PE pe33_85(.x(x85),.w(w33_84),.acc(r33_84),.res(r33_85),.clk(clk),.wout(w33_85));
	PE pe33_86(.x(x86),.w(w33_85),.acc(r33_85),.res(r33_86),.clk(clk),.wout(w33_86));
	PE pe33_87(.x(x87),.w(w33_86),.acc(r33_86),.res(r33_87),.clk(clk),.wout(w33_87));
	PE pe33_88(.x(x88),.w(w33_87),.acc(r33_87),.res(r33_88),.clk(clk),.wout(w33_88));
	PE pe33_89(.x(x89),.w(w33_88),.acc(r33_88),.res(r33_89),.clk(clk),.wout(w33_89));
	PE pe33_90(.x(x90),.w(w33_89),.acc(r33_89),.res(r33_90),.clk(clk),.wout(w33_90));
	PE pe33_91(.x(x91),.w(w33_90),.acc(r33_90),.res(r33_91),.clk(clk),.wout(w33_91));
	PE pe33_92(.x(x92),.w(w33_91),.acc(r33_91),.res(r33_92),.clk(clk),.wout(w33_92));
	PE pe33_93(.x(x93),.w(w33_92),.acc(r33_92),.res(r33_93),.clk(clk),.wout(w33_93));
	PE pe33_94(.x(x94),.w(w33_93),.acc(r33_93),.res(r33_94),.clk(clk),.wout(w33_94));
	PE pe33_95(.x(x95),.w(w33_94),.acc(r33_94),.res(r33_95),.clk(clk),.wout(w33_95));
	PE pe33_96(.x(x96),.w(w33_95),.acc(r33_95),.res(r33_96),.clk(clk),.wout(w33_96));
	PE pe33_97(.x(x97),.w(w33_96),.acc(r33_96),.res(r33_97),.clk(clk),.wout(w33_97));
	PE pe33_98(.x(x98),.w(w33_97),.acc(r33_97),.res(r33_98),.clk(clk),.wout(w33_98));
	PE pe33_99(.x(x99),.w(w33_98),.acc(r33_98),.res(r33_99),.clk(clk),.wout(w33_99));
	PE pe33_100(.x(x100),.w(w33_99),.acc(r33_99),.res(r33_100),.clk(clk),.wout(w33_100));
	PE pe33_101(.x(x101),.w(w33_100),.acc(r33_100),.res(r33_101),.clk(clk),.wout(w33_101));
	PE pe33_102(.x(x102),.w(w33_101),.acc(r33_101),.res(r33_102),.clk(clk),.wout(w33_102));
	PE pe33_103(.x(x103),.w(w33_102),.acc(r33_102),.res(r33_103),.clk(clk),.wout(w33_103));
	PE pe33_104(.x(x104),.w(w33_103),.acc(r33_103),.res(r33_104),.clk(clk),.wout(w33_104));
	PE pe33_105(.x(x105),.w(w33_104),.acc(r33_104),.res(r33_105),.clk(clk),.wout(w33_105));
	PE pe33_106(.x(x106),.w(w33_105),.acc(r33_105),.res(r33_106),.clk(clk),.wout(w33_106));
	PE pe33_107(.x(x107),.w(w33_106),.acc(r33_106),.res(r33_107),.clk(clk),.wout(w33_107));
	PE pe33_108(.x(x108),.w(w33_107),.acc(r33_107),.res(r33_108),.clk(clk),.wout(w33_108));
	PE pe33_109(.x(x109),.w(w33_108),.acc(r33_108),.res(r33_109),.clk(clk),.wout(w33_109));
	PE pe33_110(.x(x110),.w(w33_109),.acc(r33_109),.res(r33_110),.clk(clk),.wout(w33_110));
	PE pe33_111(.x(x111),.w(w33_110),.acc(r33_110),.res(r33_111),.clk(clk),.wout(w33_111));
	PE pe33_112(.x(x112),.w(w33_111),.acc(r33_111),.res(r33_112),.clk(clk),.wout(w33_112));
	PE pe33_113(.x(x113),.w(w33_112),.acc(r33_112),.res(r33_113),.clk(clk),.wout(w33_113));
	PE pe33_114(.x(x114),.w(w33_113),.acc(r33_113),.res(r33_114),.clk(clk),.wout(w33_114));
	PE pe33_115(.x(x115),.w(w33_114),.acc(r33_114),.res(r33_115),.clk(clk),.wout(w33_115));
	PE pe33_116(.x(x116),.w(w33_115),.acc(r33_115),.res(r33_116),.clk(clk),.wout(w33_116));
	PE pe33_117(.x(x117),.w(w33_116),.acc(r33_116),.res(r33_117),.clk(clk),.wout(w33_117));
	PE pe33_118(.x(x118),.w(w33_117),.acc(r33_117),.res(r33_118),.clk(clk),.wout(w33_118));
	PE pe33_119(.x(x119),.w(w33_118),.acc(r33_118),.res(r33_119),.clk(clk),.wout(w33_119));
	PE pe33_120(.x(x120),.w(w33_119),.acc(r33_119),.res(r33_120),.clk(clk),.wout(w33_120));
	PE pe33_121(.x(x121),.w(w33_120),.acc(r33_120),.res(r33_121),.clk(clk),.wout(w33_121));
	PE pe33_122(.x(x122),.w(w33_121),.acc(r33_121),.res(r33_122),.clk(clk),.wout(w33_122));
	PE pe33_123(.x(x123),.w(w33_122),.acc(r33_122),.res(r33_123),.clk(clk),.wout(w33_123));
	PE pe33_124(.x(x124),.w(w33_123),.acc(r33_123),.res(r33_124),.clk(clk),.wout(w33_124));
	PE pe33_125(.x(x125),.w(w33_124),.acc(r33_124),.res(r33_125),.clk(clk),.wout(w33_125));
	PE pe33_126(.x(x126),.w(w33_125),.acc(r33_125),.res(r33_126),.clk(clk),.wout(w33_126));
	PE pe33_127(.x(x127),.w(w33_126),.acc(r33_126),.res(result33),.clk(clk),.wout(weight33));

	PE pe34_0(.x(x0),.w(w34),.acc(32'h0),.res(r34_0),.clk(clk),.wout(w34_0));
	PE pe34_1(.x(x1),.w(w34_0),.acc(r34_0),.res(r34_1),.clk(clk),.wout(w34_1));
	PE pe34_2(.x(x2),.w(w34_1),.acc(r34_1),.res(r34_2),.clk(clk),.wout(w34_2));
	PE pe34_3(.x(x3),.w(w34_2),.acc(r34_2),.res(r34_3),.clk(clk),.wout(w34_3));
	PE pe34_4(.x(x4),.w(w34_3),.acc(r34_3),.res(r34_4),.clk(clk),.wout(w34_4));
	PE pe34_5(.x(x5),.w(w34_4),.acc(r34_4),.res(r34_5),.clk(clk),.wout(w34_5));
	PE pe34_6(.x(x6),.w(w34_5),.acc(r34_5),.res(r34_6),.clk(clk),.wout(w34_6));
	PE pe34_7(.x(x7),.w(w34_6),.acc(r34_6),.res(r34_7),.clk(clk),.wout(w34_7));
	PE pe34_8(.x(x8),.w(w34_7),.acc(r34_7),.res(r34_8),.clk(clk),.wout(w34_8));
	PE pe34_9(.x(x9),.w(w34_8),.acc(r34_8),.res(r34_9),.clk(clk),.wout(w34_9));
	PE pe34_10(.x(x10),.w(w34_9),.acc(r34_9),.res(r34_10),.clk(clk),.wout(w34_10));
	PE pe34_11(.x(x11),.w(w34_10),.acc(r34_10),.res(r34_11),.clk(clk),.wout(w34_11));
	PE pe34_12(.x(x12),.w(w34_11),.acc(r34_11),.res(r34_12),.clk(clk),.wout(w34_12));
	PE pe34_13(.x(x13),.w(w34_12),.acc(r34_12),.res(r34_13),.clk(clk),.wout(w34_13));
	PE pe34_14(.x(x14),.w(w34_13),.acc(r34_13),.res(r34_14),.clk(clk),.wout(w34_14));
	PE pe34_15(.x(x15),.w(w34_14),.acc(r34_14),.res(r34_15),.clk(clk),.wout(w34_15));
	PE pe34_16(.x(x16),.w(w34_15),.acc(r34_15),.res(r34_16),.clk(clk),.wout(w34_16));
	PE pe34_17(.x(x17),.w(w34_16),.acc(r34_16),.res(r34_17),.clk(clk),.wout(w34_17));
	PE pe34_18(.x(x18),.w(w34_17),.acc(r34_17),.res(r34_18),.clk(clk),.wout(w34_18));
	PE pe34_19(.x(x19),.w(w34_18),.acc(r34_18),.res(r34_19),.clk(clk),.wout(w34_19));
	PE pe34_20(.x(x20),.w(w34_19),.acc(r34_19),.res(r34_20),.clk(clk),.wout(w34_20));
	PE pe34_21(.x(x21),.w(w34_20),.acc(r34_20),.res(r34_21),.clk(clk),.wout(w34_21));
	PE pe34_22(.x(x22),.w(w34_21),.acc(r34_21),.res(r34_22),.clk(clk),.wout(w34_22));
	PE pe34_23(.x(x23),.w(w34_22),.acc(r34_22),.res(r34_23),.clk(clk),.wout(w34_23));
	PE pe34_24(.x(x24),.w(w34_23),.acc(r34_23),.res(r34_24),.clk(clk),.wout(w34_24));
	PE pe34_25(.x(x25),.w(w34_24),.acc(r34_24),.res(r34_25),.clk(clk),.wout(w34_25));
	PE pe34_26(.x(x26),.w(w34_25),.acc(r34_25),.res(r34_26),.clk(clk),.wout(w34_26));
	PE pe34_27(.x(x27),.w(w34_26),.acc(r34_26),.res(r34_27),.clk(clk),.wout(w34_27));
	PE pe34_28(.x(x28),.w(w34_27),.acc(r34_27),.res(r34_28),.clk(clk),.wout(w34_28));
	PE pe34_29(.x(x29),.w(w34_28),.acc(r34_28),.res(r34_29),.clk(clk),.wout(w34_29));
	PE pe34_30(.x(x30),.w(w34_29),.acc(r34_29),.res(r34_30),.clk(clk),.wout(w34_30));
	PE pe34_31(.x(x31),.w(w34_30),.acc(r34_30),.res(r34_31),.clk(clk),.wout(w34_31));
	PE pe34_32(.x(x32),.w(w34_31),.acc(r34_31),.res(r34_32),.clk(clk),.wout(w34_32));
	PE pe34_33(.x(x33),.w(w34_32),.acc(r34_32),.res(r34_33),.clk(clk),.wout(w34_33));
	PE pe34_34(.x(x34),.w(w34_33),.acc(r34_33),.res(r34_34),.clk(clk),.wout(w34_34));
	PE pe34_35(.x(x35),.w(w34_34),.acc(r34_34),.res(r34_35),.clk(clk),.wout(w34_35));
	PE pe34_36(.x(x36),.w(w34_35),.acc(r34_35),.res(r34_36),.clk(clk),.wout(w34_36));
	PE pe34_37(.x(x37),.w(w34_36),.acc(r34_36),.res(r34_37),.clk(clk),.wout(w34_37));
	PE pe34_38(.x(x38),.w(w34_37),.acc(r34_37),.res(r34_38),.clk(clk),.wout(w34_38));
	PE pe34_39(.x(x39),.w(w34_38),.acc(r34_38),.res(r34_39),.clk(clk),.wout(w34_39));
	PE pe34_40(.x(x40),.w(w34_39),.acc(r34_39),.res(r34_40),.clk(clk),.wout(w34_40));
	PE pe34_41(.x(x41),.w(w34_40),.acc(r34_40),.res(r34_41),.clk(clk),.wout(w34_41));
	PE pe34_42(.x(x42),.w(w34_41),.acc(r34_41),.res(r34_42),.clk(clk),.wout(w34_42));
	PE pe34_43(.x(x43),.w(w34_42),.acc(r34_42),.res(r34_43),.clk(clk),.wout(w34_43));
	PE pe34_44(.x(x44),.w(w34_43),.acc(r34_43),.res(r34_44),.clk(clk),.wout(w34_44));
	PE pe34_45(.x(x45),.w(w34_44),.acc(r34_44),.res(r34_45),.clk(clk),.wout(w34_45));
	PE pe34_46(.x(x46),.w(w34_45),.acc(r34_45),.res(r34_46),.clk(clk),.wout(w34_46));
	PE pe34_47(.x(x47),.w(w34_46),.acc(r34_46),.res(r34_47),.clk(clk),.wout(w34_47));
	PE pe34_48(.x(x48),.w(w34_47),.acc(r34_47),.res(r34_48),.clk(clk),.wout(w34_48));
	PE pe34_49(.x(x49),.w(w34_48),.acc(r34_48),.res(r34_49),.clk(clk),.wout(w34_49));
	PE pe34_50(.x(x50),.w(w34_49),.acc(r34_49),.res(r34_50),.clk(clk),.wout(w34_50));
	PE pe34_51(.x(x51),.w(w34_50),.acc(r34_50),.res(r34_51),.clk(clk),.wout(w34_51));
	PE pe34_52(.x(x52),.w(w34_51),.acc(r34_51),.res(r34_52),.clk(clk),.wout(w34_52));
	PE pe34_53(.x(x53),.w(w34_52),.acc(r34_52),.res(r34_53),.clk(clk),.wout(w34_53));
	PE pe34_54(.x(x54),.w(w34_53),.acc(r34_53),.res(r34_54),.clk(clk),.wout(w34_54));
	PE pe34_55(.x(x55),.w(w34_54),.acc(r34_54),.res(r34_55),.clk(clk),.wout(w34_55));
	PE pe34_56(.x(x56),.w(w34_55),.acc(r34_55),.res(r34_56),.clk(clk),.wout(w34_56));
	PE pe34_57(.x(x57),.w(w34_56),.acc(r34_56),.res(r34_57),.clk(clk),.wout(w34_57));
	PE pe34_58(.x(x58),.w(w34_57),.acc(r34_57),.res(r34_58),.clk(clk),.wout(w34_58));
	PE pe34_59(.x(x59),.w(w34_58),.acc(r34_58),.res(r34_59),.clk(clk),.wout(w34_59));
	PE pe34_60(.x(x60),.w(w34_59),.acc(r34_59),.res(r34_60),.clk(clk),.wout(w34_60));
	PE pe34_61(.x(x61),.w(w34_60),.acc(r34_60),.res(r34_61),.clk(clk),.wout(w34_61));
	PE pe34_62(.x(x62),.w(w34_61),.acc(r34_61),.res(r34_62),.clk(clk),.wout(w34_62));
	PE pe34_63(.x(x63),.w(w34_62),.acc(r34_62),.res(r34_63),.clk(clk),.wout(w34_63));
	PE pe34_64(.x(x64),.w(w34_63),.acc(r34_63),.res(r34_64),.clk(clk),.wout(w34_64));
	PE pe34_65(.x(x65),.w(w34_64),.acc(r34_64),.res(r34_65),.clk(clk),.wout(w34_65));
	PE pe34_66(.x(x66),.w(w34_65),.acc(r34_65),.res(r34_66),.clk(clk),.wout(w34_66));
	PE pe34_67(.x(x67),.w(w34_66),.acc(r34_66),.res(r34_67),.clk(clk),.wout(w34_67));
	PE pe34_68(.x(x68),.w(w34_67),.acc(r34_67),.res(r34_68),.clk(clk),.wout(w34_68));
	PE pe34_69(.x(x69),.w(w34_68),.acc(r34_68),.res(r34_69),.clk(clk),.wout(w34_69));
	PE pe34_70(.x(x70),.w(w34_69),.acc(r34_69),.res(r34_70),.clk(clk),.wout(w34_70));
	PE pe34_71(.x(x71),.w(w34_70),.acc(r34_70),.res(r34_71),.clk(clk),.wout(w34_71));
	PE pe34_72(.x(x72),.w(w34_71),.acc(r34_71),.res(r34_72),.clk(clk),.wout(w34_72));
	PE pe34_73(.x(x73),.w(w34_72),.acc(r34_72),.res(r34_73),.clk(clk),.wout(w34_73));
	PE pe34_74(.x(x74),.w(w34_73),.acc(r34_73),.res(r34_74),.clk(clk),.wout(w34_74));
	PE pe34_75(.x(x75),.w(w34_74),.acc(r34_74),.res(r34_75),.clk(clk),.wout(w34_75));
	PE pe34_76(.x(x76),.w(w34_75),.acc(r34_75),.res(r34_76),.clk(clk),.wout(w34_76));
	PE pe34_77(.x(x77),.w(w34_76),.acc(r34_76),.res(r34_77),.clk(clk),.wout(w34_77));
	PE pe34_78(.x(x78),.w(w34_77),.acc(r34_77),.res(r34_78),.clk(clk),.wout(w34_78));
	PE pe34_79(.x(x79),.w(w34_78),.acc(r34_78),.res(r34_79),.clk(clk),.wout(w34_79));
	PE pe34_80(.x(x80),.w(w34_79),.acc(r34_79),.res(r34_80),.clk(clk),.wout(w34_80));
	PE pe34_81(.x(x81),.w(w34_80),.acc(r34_80),.res(r34_81),.clk(clk),.wout(w34_81));
	PE pe34_82(.x(x82),.w(w34_81),.acc(r34_81),.res(r34_82),.clk(clk),.wout(w34_82));
	PE pe34_83(.x(x83),.w(w34_82),.acc(r34_82),.res(r34_83),.clk(clk),.wout(w34_83));
	PE pe34_84(.x(x84),.w(w34_83),.acc(r34_83),.res(r34_84),.clk(clk),.wout(w34_84));
	PE pe34_85(.x(x85),.w(w34_84),.acc(r34_84),.res(r34_85),.clk(clk),.wout(w34_85));
	PE pe34_86(.x(x86),.w(w34_85),.acc(r34_85),.res(r34_86),.clk(clk),.wout(w34_86));
	PE pe34_87(.x(x87),.w(w34_86),.acc(r34_86),.res(r34_87),.clk(clk),.wout(w34_87));
	PE pe34_88(.x(x88),.w(w34_87),.acc(r34_87),.res(r34_88),.clk(clk),.wout(w34_88));
	PE pe34_89(.x(x89),.w(w34_88),.acc(r34_88),.res(r34_89),.clk(clk),.wout(w34_89));
	PE pe34_90(.x(x90),.w(w34_89),.acc(r34_89),.res(r34_90),.clk(clk),.wout(w34_90));
	PE pe34_91(.x(x91),.w(w34_90),.acc(r34_90),.res(r34_91),.clk(clk),.wout(w34_91));
	PE pe34_92(.x(x92),.w(w34_91),.acc(r34_91),.res(r34_92),.clk(clk),.wout(w34_92));
	PE pe34_93(.x(x93),.w(w34_92),.acc(r34_92),.res(r34_93),.clk(clk),.wout(w34_93));
	PE pe34_94(.x(x94),.w(w34_93),.acc(r34_93),.res(r34_94),.clk(clk),.wout(w34_94));
	PE pe34_95(.x(x95),.w(w34_94),.acc(r34_94),.res(r34_95),.clk(clk),.wout(w34_95));
	PE pe34_96(.x(x96),.w(w34_95),.acc(r34_95),.res(r34_96),.clk(clk),.wout(w34_96));
	PE pe34_97(.x(x97),.w(w34_96),.acc(r34_96),.res(r34_97),.clk(clk),.wout(w34_97));
	PE pe34_98(.x(x98),.w(w34_97),.acc(r34_97),.res(r34_98),.clk(clk),.wout(w34_98));
	PE pe34_99(.x(x99),.w(w34_98),.acc(r34_98),.res(r34_99),.clk(clk),.wout(w34_99));
	PE pe34_100(.x(x100),.w(w34_99),.acc(r34_99),.res(r34_100),.clk(clk),.wout(w34_100));
	PE pe34_101(.x(x101),.w(w34_100),.acc(r34_100),.res(r34_101),.clk(clk),.wout(w34_101));
	PE pe34_102(.x(x102),.w(w34_101),.acc(r34_101),.res(r34_102),.clk(clk),.wout(w34_102));
	PE pe34_103(.x(x103),.w(w34_102),.acc(r34_102),.res(r34_103),.clk(clk),.wout(w34_103));
	PE pe34_104(.x(x104),.w(w34_103),.acc(r34_103),.res(r34_104),.clk(clk),.wout(w34_104));
	PE pe34_105(.x(x105),.w(w34_104),.acc(r34_104),.res(r34_105),.clk(clk),.wout(w34_105));
	PE pe34_106(.x(x106),.w(w34_105),.acc(r34_105),.res(r34_106),.clk(clk),.wout(w34_106));
	PE pe34_107(.x(x107),.w(w34_106),.acc(r34_106),.res(r34_107),.clk(clk),.wout(w34_107));
	PE pe34_108(.x(x108),.w(w34_107),.acc(r34_107),.res(r34_108),.clk(clk),.wout(w34_108));
	PE pe34_109(.x(x109),.w(w34_108),.acc(r34_108),.res(r34_109),.clk(clk),.wout(w34_109));
	PE pe34_110(.x(x110),.w(w34_109),.acc(r34_109),.res(r34_110),.clk(clk),.wout(w34_110));
	PE pe34_111(.x(x111),.w(w34_110),.acc(r34_110),.res(r34_111),.clk(clk),.wout(w34_111));
	PE pe34_112(.x(x112),.w(w34_111),.acc(r34_111),.res(r34_112),.clk(clk),.wout(w34_112));
	PE pe34_113(.x(x113),.w(w34_112),.acc(r34_112),.res(r34_113),.clk(clk),.wout(w34_113));
	PE pe34_114(.x(x114),.w(w34_113),.acc(r34_113),.res(r34_114),.clk(clk),.wout(w34_114));
	PE pe34_115(.x(x115),.w(w34_114),.acc(r34_114),.res(r34_115),.clk(clk),.wout(w34_115));
	PE pe34_116(.x(x116),.w(w34_115),.acc(r34_115),.res(r34_116),.clk(clk),.wout(w34_116));
	PE pe34_117(.x(x117),.w(w34_116),.acc(r34_116),.res(r34_117),.clk(clk),.wout(w34_117));
	PE pe34_118(.x(x118),.w(w34_117),.acc(r34_117),.res(r34_118),.clk(clk),.wout(w34_118));
	PE pe34_119(.x(x119),.w(w34_118),.acc(r34_118),.res(r34_119),.clk(clk),.wout(w34_119));
	PE pe34_120(.x(x120),.w(w34_119),.acc(r34_119),.res(r34_120),.clk(clk),.wout(w34_120));
	PE pe34_121(.x(x121),.w(w34_120),.acc(r34_120),.res(r34_121),.clk(clk),.wout(w34_121));
	PE pe34_122(.x(x122),.w(w34_121),.acc(r34_121),.res(r34_122),.clk(clk),.wout(w34_122));
	PE pe34_123(.x(x123),.w(w34_122),.acc(r34_122),.res(r34_123),.clk(clk),.wout(w34_123));
	PE pe34_124(.x(x124),.w(w34_123),.acc(r34_123),.res(r34_124),.clk(clk),.wout(w34_124));
	PE pe34_125(.x(x125),.w(w34_124),.acc(r34_124),.res(r34_125),.clk(clk),.wout(w34_125));
	PE pe34_126(.x(x126),.w(w34_125),.acc(r34_125),.res(r34_126),.clk(clk),.wout(w34_126));
	PE pe34_127(.x(x127),.w(w34_126),.acc(r34_126),.res(result34),.clk(clk),.wout(weight34));

	PE pe35_0(.x(x0),.w(w35),.acc(32'h0),.res(r35_0),.clk(clk),.wout(w35_0));
	PE pe35_1(.x(x1),.w(w35_0),.acc(r35_0),.res(r35_1),.clk(clk),.wout(w35_1));
	PE pe35_2(.x(x2),.w(w35_1),.acc(r35_1),.res(r35_2),.clk(clk),.wout(w35_2));
	PE pe35_3(.x(x3),.w(w35_2),.acc(r35_2),.res(r35_3),.clk(clk),.wout(w35_3));
	PE pe35_4(.x(x4),.w(w35_3),.acc(r35_3),.res(r35_4),.clk(clk),.wout(w35_4));
	PE pe35_5(.x(x5),.w(w35_4),.acc(r35_4),.res(r35_5),.clk(clk),.wout(w35_5));
	PE pe35_6(.x(x6),.w(w35_5),.acc(r35_5),.res(r35_6),.clk(clk),.wout(w35_6));
	PE pe35_7(.x(x7),.w(w35_6),.acc(r35_6),.res(r35_7),.clk(clk),.wout(w35_7));
	PE pe35_8(.x(x8),.w(w35_7),.acc(r35_7),.res(r35_8),.clk(clk),.wout(w35_8));
	PE pe35_9(.x(x9),.w(w35_8),.acc(r35_8),.res(r35_9),.clk(clk),.wout(w35_9));
	PE pe35_10(.x(x10),.w(w35_9),.acc(r35_9),.res(r35_10),.clk(clk),.wout(w35_10));
	PE pe35_11(.x(x11),.w(w35_10),.acc(r35_10),.res(r35_11),.clk(clk),.wout(w35_11));
	PE pe35_12(.x(x12),.w(w35_11),.acc(r35_11),.res(r35_12),.clk(clk),.wout(w35_12));
	PE pe35_13(.x(x13),.w(w35_12),.acc(r35_12),.res(r35_13),.clk(clk),.wout(w35_13));
	PE pe35_14(.x(x14),.w(w35_13),.acc(r35_13),.res(r35_14),.clk(clk),.wout(w35_14));
	PE pe35_15(.x(x15),.w(w35_14),.acc(r35_14),.res(r35_15),.clk(clk),.wout(w35_15));
	PE pe35_16(.x(x16),.w(w35_15),.acc(r35_15),.res(r35_16),.clk(clk),.wout(w35_16));
	PE pe35_17(.x(x17),.w(w35_16),.acc(r35_16),.res(r35_17),.clk(clk),.wout(w35_17));
	PE pe35_18(.x(x18),.w(w35_17),.acc(r35_17),.res(r35_18),.clk(clk),.wout(w35_18));
	PE pe35_19(.x(x19),.w(w35_18),.acc(r35_18),.res(r35_19),.clk(clk),.wout(w35_19));
	PE pe35_20(.x(x20),.w(w35_19),.acc(r35_19),.res(r35_20),.clk(clk),.wout(w35_20));
	PE pe35_21(.x(x21),.w(w35_20),.acc(r35_20),.res(r35_21),.clk(clk),.wout(w35_21));
	PE pe35_22(.x(x22),.w(w35_21),.acc(r35_21),.res(r35_22),.clk(clk),.wout(w35_22));
	PE pe35_23(.x(x23),.w(w35_22),.acc(r35_22),.res(r35_23),.clk(clk),.wout(w35_23));
	PE pe35_24(.x(x24),.w(w35_23),.acc(r35_23),.res(r35_24),.clk(clk),.wout(w35_24));
	PE pe35_25(.x(x25),.w(w35_24),.acc(r35_24),.res(r35_25),.clk(clk),.wout(w35_25));
	PE pe35_26(.x(x26),.w(w35_25),.acc(r35_25),.res(r35_26),.clk(clk),.wout(w35_26));
	PE pe35_27(.x(x27),.w(w35_26),.acc(r35_26),.res(r35_27),.clk(clk),.wout(w35_27));
	PE pe35_28(.x(x28),.w(w35_27),.acc(r35_27),.res(r35_28),.clk(clk),.wout(w35_28));
	PE pe35_29(.x(x29),.w(w35_28),.acc(r35_28),.res(r35_29),.clk(clk),.wout(w35_29));
	PE pe35_30(.x(x30),.w(w35_29),.acc(r35_29),.res(r35_30),.clk(clk),.wout(w35_30));
	PE pe35_31(.x(x31),.w(w35_30),.acc(r35_30),.res(r35_31),.clk(clk),.wout(w35_31));
	PE pe35_32(.x(x32),.w(w35_31),.acc(r35_31),.res(r35_32),.clk(clk),.wout(w35_32));
	PE pe35_33(.x(x33),.w(w35_32),.acc(r35_32),.res(r35_33),.clk(clk),.wout(w35_33));
	PE pe35_34(.x(x34),.w(w35_33),.acc(r35_33),.res(r35_34),.clk(clk),.wout(w35_34));
	PE pe35_35(.x(x35),.w(w35_34),.acc(r35_34),.res(r35_35),.clk(clk),.wout(w35_35));
	PE pe35_36(.x(x36),.w(w35_35),.acc(r35_35),.res(r35_36),.clk(clk),.wout(w35_36));
	PE pe35_37(.x(x37),.w(w35_36),.acc(r35_36),.res(r35_37),.clk(clk),.wout(w35_37));
	PE pe35_38(.x(x38),.w(w35_37),.acc(r35_37),.res(r35_38),.clk(clk),.wout(w35_38));
	PE pe35_39(.x(x39),.w(w35_38),.acc(r35_38),.res(r35_39),.clk(clk),.wout(w35_39));
	PE pe35_40(.x(x40),.w(w35_39),.acc(r35_39),.res(r35_40),.clk(clk),.wout(w35_40));
	PE pe35_41(.x(x41),.w(w35_40),.acc(r35_40),.res(r35_41),.clk(clk),.wout(w35_41));
	PE pe35_42(.x(x42),.w(w35_41),.acc(r35_41),.res(r35_42),.clk(clk),.wout(w35_42));
	PE pe35_43(.x(x43),.w(w35_42),.acc(r35_42),.res(r35_43),.clk(clk),.wout(w35_43));
	PE pe35_44(.x(x44),.w(w35_43),.acc(r35_43),.res(r35_44),.clk(clk),.wout(w35_44));
	PE pe35_45(.x(x45),.w(w35_44),.acc(r35_44),.res(r35_45),.clk(clk),.wout(w35_45));
	PE pe35_46(.x(x46),.w(w35_45),.acc(r35_45),.res(r35_46),.clk(clk),.wout(w35_46));
	PE pe35_47(.x(x47),.w(w35_46),.acc(r35_46),.res(r35_47),.clk(clk),.wout(w35_47));
	PE pe35_48(.x(x48),.w(w35_47),.acc(r35_47),.res(r35_48),.clk(clk),.wout(w35_48));
	PE pe35_49(.x(x49),.w(w35_48),.acc(r35_48),.res(r35_49),.clk(clk),.wout(w35_49));
	PE pe35_50(.x(x50),.w(w35_49),.acc(r35_49),.res(r35_50),.clk(clk),.wout(w35_50));
	PE pe35_51(.x(x51),.w(w35_50),.acc(r35_50),.res(r35_51),.clk(clk),.wout(w35_51));
	PE pe35_52(.x(x52),.w(w35_51),.acc(r35_51),.res(r35_52),.clk(clk),.wout(w35_52));
	PE pe35_53(.x(x53),.w(w35_52),.acc(r35_52),.res(r35_53),.clk(clk),.wout(w35_53));
	PE pe35_54(.x(x54),.w(w35_53),.acc(r35_53),.res(r35_54),.clk(clk),.wout(w35_54));
	PE pe35_55(.x(x55),.w(w35_54),.acc(r35_54),.res(r35_55),.clk(clk),.wout(w35_55));
	PE pe35_56(.x(x56),.w(w35_55),.acc(r35_55),.res(r35_56),.clk(clk),.wout(w35_56));
	PE pe35_57(.x(x57),.w(w35_56),.acc(r35_56),.res(r35_57),.clk(clk),.wout(w35_57));
	PE pe35_58(.x(x58),.w(w35_57),.acc(r35_57),.res(r35_58),.clk(clk),.wout(w35_58));
	PE pe35_59(.x(x59),.w(w35_58),.acc(r35_58),.res(r35_59),.clk(clk),.wout(w35_59));
	PE pe35_60(.x(x60),.w(w35_59),.acc(r35_59),.res(r35_60),.clk(clk),.wout(w35_60));
	PE pe35_61(.x(x61),.w(w35_60),.acc(r35_60),.res(r35_61),.clk(clk),.wout(w35_61));
	PE pe35_62(.x(x62),.w(w35_61),.acc(r35_61),.res(r35_62),.clk(clk),.wout(w35_62));
	PE pe35_63(.x(x63),.w(w35_62),.acc(r35_62),.res(r35_63),.clk(clk),.wout(w35_63));
	PE pe35_64(.x(x64),.w(w35_63),.acc(r35_63),.res(r35_64),.clk(clk),.wout(w35_64));
	PE pe35_65(.x(x65),.w(w35_64),.acc(r35_64),.res(r35_65),.clk(clk),.wout(w35_65));
	PE pe35_66(.x(x66),.w(w35_65),.acc(r35_65),.res(r35_66),.clk(clk),.wout(w35_66));
	PE pe35_67(.x(x67),.w(w35_66),.acc(r35_66),.res(r35_67),.clk(clk),.wout(w35_67));
	PE pe35_68(.x(x68),.w(w35_67),.acc(r35_67),.res(r35_68),.clk(clk),.wout(w35_68));
	PE pe35_69(.x(x69),.w(w35_68),.acc(r35_68),.res(r35_69),.clk(clk),.wout(w35_69));
	PE pe35_70(.x(x70),.w(w35_69),.acc(r35_69),.res(r35_70),.clk(clk),.wout(w35_70));
	PE pe35_71(.x(x71),.w(w35_70),.acc(r35_70),.res(r35_71),.clk(clk),.wout(w35_71));
	PE pe35_72(.x(x72),.w(w35_71),.acc(r35_71),.res(r35_72),.clk(clk),.wout(w35_72));
	PE pe35_73(.x(x73),.w(w35_72),.acc(r35_72),.res(r35_73),.clk(clk),.wout(w35_73));
	PE pe35_74(.x(x74),.w(w35_73),.acc(r35_73),.res(r35_74),.clk(clk),.wout(w35_74));
	PE pe35_75(.x(x75),.w(w35_74),.acc(r35_74),.res(r35_75),.clk(clk),.wout(w35_75));
	PE pe35_76(.x(x76),.w(w35_75),.acc(r35_75),.res(r35_76),.clk(clk),.wout(w35_76));
	PE pe35_77(.x(x77),.w(w35_76),.acc(r35_76),.res(r35_77),.clk(clk),.wout(w35_77));
	PE pe35_78(.x(x78),.w(w35_77),.acc(r35_77),.res(r35_78),.clk(clk),.wout(w35_78));
	PE pe35_79(.x(x79),.w(w35_78),.acc(r35_78),.res(r35_79),.clk(clk),.wout(w35_79));
	PE pe35_80(.x(x80),.w(w35_79),.acc(r35_79),.res(r35_80),.clk(clk),.wout(w35_80));
	PE pe35_81(.x(x81),.w(w35_80),.acc(r35_80),.res(r35_81),.clk(clk),.wout(w35_81));
	PE pe35_82(.x(x82),.w(w35_81),.acc(r35_81),.res(r35_82),.clk(clk),.wout(w35_82));
	PE pe35_83(.x(x83),.w(w35_82),.acc(r35_82),.res(r35_83),.clk(clk),.wout(w35_83));
	PE pe35_84(.x(x84),.w(w35_83),.acc(r35_83),.res(r35_84),.clk(clk),.wout(w35_84));
	PE pe35_85(.x(x85),.w(w35_84),.acc(r35_84),.res(r35_85),.clk(clk),.wout(w35_85));
	PE pe35_86(.x(x86),.w(w35_85),.acc(r35_85),.res(r35_86),.clk(clk),.wout(w35_86));
	PE pe35_87(.x(x87),.w(w35_86),.acc(r35_86),.res(r35_87),.clk(clk),.wout(w35_87));
	PE pe35_88(.x(x88),.w(w35_87),.acc(r35_87),.res(r35_88),.clk(clk),.wout(w35_88));
	PE pe35_89(.x(x89),.w(w35_88),.acc(r35_88),.res(r35_89),.clk(clk),.wout(w35_89));
	PE pe35_90(.x(x90),.w(w35_89),.acc(r35_89),.res(r35_90),.clk(clk),.wout(w35_90));
	PE pe35_91(.x(x91),.w(w35_90),.acc(r35_90),.res(r35_91),.clk(clk),.wout(w35_91));
	PE pe35_92(.x(x92),.w(w35_91),.acc(r35_91),.res(r35_92),.clk(clk),.wout(w35_92));
	PE pe35_93(.x(x93),.w(w35_92),.acc(r35_92),.res(r35_93),.clk(clk),.wout(w35_93));
	PE pe35_94(.x(x94),.w(w35_93),.acc(r35_93),.res(r35_94),.clk(clk),.wout(w35_94));
	PE pe35_95(.x(x95),.w(w35_94),.acc(r35_94),.res(r35_95),.clk(clk),.wout(w35_95));
	PE pe35_96(.x(x96),.w(w35_95),.acc(r35_95),.res(r35_96),.clk(clk),.wout(w35_96));
	PE pe35_97(.x(x97),.w(w35_96),.acc(r35_96),.res(r35_97),.clk(clk),.wout(w35_97));
	PE pe35_98(.x(x98),.w(w35_97),.acc(r35_97),.res(r35_98),.clk(clk),.wout(w35_98));
	PE pe35_99(.x(x99),.w(w35_98),.acc(r35_98),.res(r35_99),.clk(clk),.wout(w35_99));
	PE pe35_100(.x(x100),.w(w35_99),.acc(r35_99),.res(r35_100),.clk(clk),.wout(w35_100));
	PE pe35_101(.x(x101),.w(w35_100),.acc(r35_100),.res(r35_101),.clk(clk),.wout(w35_101));
	PE pe35_102(.x(x102),.w(w35_101),.acc(r35_101),.res(r35_102),.clk(clk),.wout(w35_102));
	PE pe35_103(.x(x103),.w(w35_102),.acc(r35_102),.res(r35_103),.clk(clk),.wout(w35_103));
	PE pe35_104(.x(x104),.w(w35_103),.acc(r35_103),.res(r35_104),.clk(clk),.wout(w35_104));
	PE pe35_105(.x(x105),.w(w35_104),.acc(r35_104),.res(r35_105),.clk(clk),.wout(w35_105));
	PE pe35_106(.x(x106),.w(w35_105),.acc(r35_105),.res(r35_106),.clk(clk),.wout(w35_106));
	PE pe35_107(.x(x107),.w(w35_106),.acc(r35_106),.res(r35_107),.clk(clk),.wout(w35_107));
	PE pe35_108(.x(x108),.w(w35_107),.acc(r35_107),.res(r35_108),.clk(clk),.wout(w35_108));
	PE pe35_109(.x(x109),.w(w35_108),.acc(r35_108),.res(r35_109),.clk(clk),.wout(w35_109));
	PE pe35_110(.x(x110),.w(w35_109),.acc(r35_109),.res(r35_110),.clk(clk),.wout(w35_110));
	PE pe35_111(.x(x111),.w(w35_110),.acc(r35_110),.res(r35_111),.clk(clk),.wout(w35_111));
	PE pe35_112(.x(x112),.w(w35_111),.acc(r35_111),.res(r35_112),.clk(clk),.wout(w35_112));
	PE pe35_113(.x(x113),.w(w35_112),.acc(r35_112),.res(r35_113),.clk(clk),.wout(w35_113));
	PE pe35_114(.x(x114),.w(w35_113),.acc(r35_113),.res(r35_114),.clk(clk),.wout(w35_114));
	PE pe35_115(.x(x115),.w(w35_114),.acc(r35_114),.res(r35_115),.clk(clk),.wout(w35_115));
	PE pe35_116(.x(x116),.w(w35_115),.acc(r35_115),.res(r35_116),.clk(clk),.wout(w35_116));
	PE pe35_117(.x(x117),.w(w35_116),.acc(r35_116),.res(r35_117),.clk(clk),.wout(w35_117));
	PE pe35_118(.x(x118),.w(w35_117),.acc(r35_117),.res(r35_118),.clk(clk),.wout(w35_118));
	PE pe35_119(.x(x119),.w(w35_118),.acc(r35_118),.res(r35_119),.clk(clk),.wout(w35_119));
	PE pe35_120(.x(x120),.w(w35_119),.acc(r35_119),.res(r35_120),.clk(clk),.wout(w35_120));
	PE pe35_121(.x(x121),.w(w35_120),.acc(r35_120),.res(r35_121),.clk(clk),.wout(w35_121));
	PE pe35_122(.x(x122),.w(w35_121),.acc(r35_121),.res(r35_122),.clk(clk),.wout(w35_122));
	PE pe35_123(.x(x123),.w(w35_122),.acc(r35_122),.res(r35_123),.clk(clk),.wout(w35_123));
	PE pe35_124(.x(x124),.w(w35_123),.acc(r35_123),.res(r35_124),.clk(clk),.wout(w35_124));
	PE pe35_125(.x(x125),.w(w35_124),.acc(r35_124),.res(r35_125),.clk(clk),.wout(w35_125));
	PE pe35_126(.x(x126),.w(w35_125),.acc(r35_125),.res(r35_126),.clk(clk),.wout(w35_126));
	PE pe35_127(.x(x127),.w(w35_126),.acc(r35_126),.res(result35),.clk(clk),.wout(weight35));

	PE pe36_0(.x(x0),.w(w36),.acc(32'h0),.res(r36_0),.clk(clk),.wout(w36_0));
	PE pe36_1(.x(x1),.w(w36_0),.acc(r36_0),.res(r36_1),.clk(clk),.wout(w36_1));
	PE pe36_2(.x(x2),.w(w36_1),.acc(r36_1),.res(r36_2),.clk(clk),.wout(w36_2));
	PE pe36_3(.x(x3),.w(w36_2),.acc(r36_2),.res(r36_3),.clk(clk),.wout(w36_3));
	PE pe36_4(.x(x4),.w(w36_3),.acc(r36_3),.res(r36_4),.clk(clk),.wout(w36_4));
	PE pe36_5(.x(x5),.w(w36_4),.acc(r36_4),.res(r36_5),.clk(clk),.wout(w36_5));
	PE pe36_6(.x(x6),.w(w36_5),.acc(r36_5),.res(r36_6),.clk(clk),.wout(w36_6));
	PE pe36_7(.x(x7),.w(w36_6),.acc(r36_6),.res(r36_7),.clk(clk),.wout(w36_7));
	PE pe36_8(.x(x8),.w(w36_7),.acc(r36_7),.res(r36_8),.clk(clk),.wout(w36_8));
	PE pe36_9(.x(x9),.w(w36_8),.acc(r36_8),.res(r36_9),.clk(clk),.wout(w36_9));
	PE pe36_10(.x(x10),.w(w36_9),.acc(r36_9),.res(r36_10),.clk(clk),.wout(w36_10));
	PE pe36_11(.x(x11),.w(w36_10),.acc(r36_10),.res(r36_11),.clk(clk),.wout(w36_11));
	PE pe36_12(.x(x12),.w(w36_11),.acc(r36_11),.res(r36_12),.clk(clk),.wout(w36_12));
	PE pe36_13(.x(x13),.w(w36_12),.acc(r36_12),.res(r36_13),.clk(clk),.wout(w36_13));
	PE pe36_14(.x(x14),.w(w36_13),.acc(r36_13),.res(r36_14),.clk(clk),.wout(w36_14));
	PE pe36_15(.x(x15),.w(w36_14),.acc(r36_14),.res(r36_15),.clk(clk),.wout(w36_15));
	PE pe36_16(.x(x16),.w(w36_15),.acc(r36_15),.res(r36_16),.clk(clk),.wout(w36_16));
	PE pe36_17(.x(x17),.w(w36_16),.acc(r36_16),.res(r36_17),.clk(clk),.wout(w36_17));
	PE pe36_18(.x(x18),.w(w36_17),.acc(r36_17),.res(r36_18),.clk(clk),.wout(w36_18));
	PE pe36_19(.x(x19),.w(w36_18),.acc(r36_18),.res(r36_19),.clk(clk),.wout(w36_19));
	PE pe36_20(.x(x20),.w(w36_19),.acc(r36_19),.res(r36_20),.clk(clk),.wout(w36_20));
	PE pe36_21(.x(x21),.w(w36_20),.acc(r36_20),.res(r36_21),.clk(clk),.wout(w36_21));
	PE pe36_22(.x(x22),.w(w36_21),.acc(r36_21),.res(r36_22),.clk(clk),.wout(w36_22));
	PE pe36_23(.x(x23),.w(w36_22),.acc(r36_22),.res(r36_23),.clk(clk),.wout(w36_23));
	PE pe36_24(.x(x24),.w(w36_23),.acc(r36_23),.res(r36_24),.clk(clk),.wout(w36_24));
	PE pe36_25(.x(x25),.w(w36_24),.acc(r36_24),.res(r36_25),.clk(clk),.wout(w36_25));
	PE pe36_26(.x(x26),.w(w36_25),.acc(r36_25),.res(r36_26),.clk(clk),.wout(w36_26));
	PE pe36_27(.x(x27),.w(w36_26),.acc(r36_26),.res(r36_27),.clk(clk),.wout(w36_27));
	PE pe36_28(.x(x28),.w(w36_27),.acc(r36_27),.res(r36_28),.clk(clk),.wout(w36_28));
	PE pe36_29(.x(x29),.w(w36_28),.acc(r36_28),.res(r36_29),.clk(clk),.wout(w36_29));
	PE pe36_30(.x(x30),.w(w36_29),.acc(r36_29),.res(r36_30),.clk(clk),.wout(w36_30));
	PE pe36_31(.x(x31),.w(w36_30),.acc(r36_30),.res(r36_31),.clk(clk),.wout(w36_31));
	PE pe36_32(.x(x32),.w(w36_31),.acc(r36_31),.res(r36_32),.clk(clk),.wout(w36_32));
	PE pe36_33(.x(x33),.w(w36_32),.acc(r36_32),.res(r36_33),.clk(clk),.wout(w36_33));
	PE pe36_34(.x(x34),.w(w36_33),.acc(r36_33),.res(r36_34),.clk(clk),.wout(w36_34));
	PE pe36_35(.x(x35),.w(w36_34),.acc(r36_34),.res(r36_35),.clk(clk),.wout(w36_35));
	PE pe36_36(.x(x36),.w(w36_35),.acc(r36_35),.res(r36_36),.clk(clk),.wout(w36_36));
	PE pe36_37(.x(x37),.w(w36_36),.acc(r36_36),.res(r36_37),.clk(clk),.wout(w36_37));
	PE pe36_38(.x(x38),.w(w36_37),.acc(r36_37),.res(r36_38),.clk(clk),.wout(w36_38));
	PE pe36_39(.x(x39),.w(w36_38),.acc(r36_38),.res(r36_39),.clk(clk),.wout(w36_39));
	PE pe36_40(.x(x40),.w(w36_39),.acc(r36_39),.res(r36_40),.clk(clk),.wout(w36_40));
	PE pe36_41(.x(x41),.w(w36_40),.acc(r36_40),.res(r36_41),.clk(clk),.wout(w36_41));
	PE pe36_42(.x(x42),.w(w36_41),.acc(r36_41),.res(r36_42),.clk(clk),.wout(w36_42));
	PE pe36_43(.x(x43),.w(w36_42),.acc(r36_42),.res(r36_43),.clk(clk),.wout(w36_43));
	PE pe36_44(.x(x44),.w(w36_43),.acc(r36_43),.res(r36_44),.clk(clk),.wout(w36_44));
	PE pe36_45(.x(x45),.w(w36_44),.acc(r36_44),.res(r36_45),.clk(clk),.wout(w36_45));
	PE pe36_46(.x(x46),.w(w36_45),.acc(r36_45),.res(r36_46),.clk(clk),.wout(w36_46));
	PE pe36_47(.x(x47),.w(w36_46),.acc(r36_46),.res(r36_47),.clk(clk),.wout(w36_47));
	PE pe36_48(.x(x48),.w(w36_47),.acc(r36_47),.res(r36_48),.clk(clk),.wout(w36_48));
	PE pe36_49(.x(x49),.w(w36_48),.acc(r36_48),.res(r36_49),.clk(clk),.wout(w36_49));
	PE pe36_50(.x(x50),.w(w36_49),.acc(r36_49),.res(r36_50),.clk(clk),.wout(w36_50));
	PE pe36_51(.x(x51),.w(w36_50),.acc(r36_50),.res(r36_51),.clk(clk),.wout(w36_51));
	PE pe36_52(.x(x52),.w(w36_51),.acc(r36_51),.res(r36_52),.clk(clk),.wout(w36_52));
	PE pe36_53(.x(x53),.w(w36_52),.acc(r36_52),.res(r36_53),.clk(clk),.wout(w36_53));
	PE pe36_54(.x(x54),.w(w36_53),.acc(r36_53),.res(r36_54),.clk(clk),.wout(w36_54));
	PE pe36_55(.x(x55),.w(w36_54),.acc(r36_54),.res(r36_55),.clk(clk),.wout(w36_55));
	PE pe36_56(.x(x56),.w(w36_55),.acc(r36_55),.res(r36_56),.clk(clk),.wout(w36_56));
	PE pe36_57(.x(x57),.w(w36_56),.acc(r36_56),.res(r36_57),.clk(clk),.wout(w36_57));
	PE pe36_58(.x(x58),.w(w36_57),.acc(r36_57),.res(r36_58),.clk(clk),.wout(w36_58));
	PE pe36_59(.x(x59),.w(w36_58),.acc(r36_58),.res(r36_59),.clk(clk),.wout(w36_59));
	PE pe36_60(.x(x60),.w(w36_59),.acc(r36_59),.res(r36_60),.clk(clk),.wout(w36_60));
	PE pe36_61(.x(x61),.w(w36_60),.acc(r36_60),.res(r36_61),.clk(clk),.wout(w36_61));
	PE pe36_62(.x(x62),.w(w36_61),.acc(r36_61),.res(r36_62),.clk(clk),.wout(w36_62));
	PE pe36_63(.x(x63),.w(w36_62),.acc(r36_62),.res(r36_63),.clk(clk),.wout(w36_63));
	PE pe36_64(.x(x64),.w(w36_63),.acc(r36_63),.res(r36_64),.clk(clk),.wout(w36_64));
	PE pe36_65(.x(x65),.w(w36_64),.acc(r36_64),.res(r36_65),.clk(clk),.wout(w36_65));
	PE pe36_66(.x(x66),.w(w36_65),.acc(r36_65),.res(r36_66),.clk(clk),.wout(w36_66));
	PE pe36_67(.x(x67),.w(w36_66),.acc(r36_66),.res(r36_67),.clk(clk),.wout(w36_67));
	PE pe36_68(.x(x68),.w(w36_67),.acc(r36_67),.res(r36_68),.clk(clk),.wout(w36_68));
	PE pe36_69(.x(x69),.w(w36_68),.acc(r36_68),.res(r36_69),.clk(clk),.wout(w36_69));
	PE pe36_70(.x(x70),.w(w36_69),.acc(r36_69),.res(r36_70),.clk(clk),.wout(w36_70));
	PE pe36_71(.x(x71),.w(w36_70),.acc(r36_70),.res(r36_71),.clk(clk),.wout(w36_71));
	PE pe36_72(.x(x72),.w(w36_71),.acc(r36_71),.res(r36_72),.clk(clk),.wout(w36_72));
	PE pe36_73(.x(x73),.w(w36_72),.acc(r36_72),.res(r36_73),.clk(clk),.wout(w36_73));
	PE pe36_74(.x(x74),.w(w36_73),.acc(r36_73),.res(r36_74),.clk(clk),.wout(w36_74));
	PE pe36_75(.x(x75),.w(w36_74),.acc(r36_74),.res(r36_75),.clk(clk),.wout(w36_75));
	PE pe36_76(.x(x76),.w(w36_75),.acc(r36_75),.res(r36_76),.clk(clk),.wout(w36_76));
	PE pe36_77(.x(x77),.w(w36_76),.acc(r36_76),.res(r36_77),.clk(clk),.wout(w36_77));
	PE pe36_78(.x(x78),.w(w36_77),.acc(r36_77),.res(r36_78),.clk(clk),.wout(w36_78));
	PE pe36_79(.x(x79),.w(w36_78),.acc(r36_78),.res(r36_79),.clk(clk),.wout(w36_79));
	PE pe36_80(.x(x80),.w(w36_79),.acc(r36_79),.res(r36_80),.clk(clk),.wout(w36_80));
	PE pe36_81(.x(x81),.w(w36_80),.acc(r36_80),.res(r36_81),.clk(clk),.wout(w36_81));
	PE pe36_82(.x(x82),.w(w36_81),.acc(r36_81),.res(r36_82),.clk(clk),.wout(w36_82));
	PE pe36_83(.x(x83),.w(w36_82),.acc(r36_82),.res(r36_83),.clk(clk),.wout(w36_83));
	PE pe36_84(.x(x84),.w(w36_83),.acc(r36_83),.res(r36_84),.clk(clk),.wout(w36_84));
	PE pe36_85(.x(x85),.w(w36_84),.acc(r36_84),.res(r36_85),.clk(clk),.wout(w36_85));
	PE pe36_86(.x(x86),.w(w36_85),.acc(r36_85),.res(r36_86),.clk(clk),.wout(w36_86));
	PE pe36_87(.x(x87),.w(w36_86),.acc(r36_86),.res(r36_87),.clk(clk),.wout(w36_87));
	PE pe36_88(.x(x88),.w(w36_87),.acc(r36_87),.res(r36_88),.clk(clk),.wout(w36_88));
	PE pe36_89(.x(x89),.w(w36_88),.acc(r36_88),.res(r36_89),.clk(clk),.wout(w36_89));
	PE pe36_90(.x(x90),.w(w36_89),.acc(r36_89),.res(r36_90),.clk(clk),.wout(w36_90));
	PE pe36_91(.x(x91),.w(w36_90),.acc(r36_90),.res(r36_91),.clk(clk),.wout(w36_91));
	PE pe36_92(.x(x92),.w(w36_91),.acc(r36_91),.res(r36_92),.clk(clk),.wout(w36_92));
	PE pe36_93(.x(x93),.w(w36_92),.acc(r36_92),.res(r36_93),.clk(clk),.wout(w36_93));
	PE pe36_94(.x(x94),.w(w36_93),.acc(r36_93),.res(r36_94),.clk(clk),.wout(w36_94));
	PE pe36_95(.x(x95),.w(w36_94),.acc(r36_94),.res(r36_95),.clk(clk),.wout(w36_95));
	PE pe36_96(.x(x96),.w(w36_95),.acc(r36_95),.res(r36_96),.clk(clk),.wout(w36_96));
	PE pe36_97(.x(x97),.w(w36_96),.acc(r36_96),.res(r36_97),.clk(clk),.wout(w36_97));
	PE pe36_98(.x(x98),.w(w36_97),.acc(r36_97),.res(r36_98),.clk(clk),.wout(w36_98));
	PE pe36_99(.x(x99),.w(w36_98),.acc(r36_98),.res(r36_99),.clk(clk),.wout(w36_99));
	PE pe36_100(.x(x100),.w(w36_99),.acc(r36_99),.res(r36_100),.clk(clk),.wout(w36_100));
	PE pe36_101(.x(x101),.w(w36_100),.acc(r36_100),.res(r36_101),.clk(clk),.wout(w36_101));
	PE pe36_102(.x(x102),.w(w36_101),.acc(r36_101),.res(r36_102),.clk(clk),.wout(w36_102));
	PE pe36_103(.x(x103),.w(w36_102),.acc(r36_102),.res(r36_103),.clk(clk),.wout(w36_103));
	PE pe36_104(.x(x104),.w(w36_103),.acc(r36_103),.res(r36_104),.clk(clk),.wout(w36_104));
	PE pe36_105(.x(x105),.w(w36_104),.acc(r36_104),.res(r36_105),.clk(clk),.wout(w36_105));
	PE pe36_106(.x(x106),.w(w36_105),.acc(r36_105),.res(r36_106),.clk(clk),.wout(w36_106));
	PE pe36_107(.x(x107),.w(w36_106),.acc(r36_106),.res(r36_107),.clk(clk),.wout(w36_107));
	PE pe36_108(.x(x108),.w(w36_107),.acc(r36_107),.res(r36_108),.clk(clk),.wout(w36_108));
	PE pe36_109(.x(x109),.w(w36_108),.acc(r36_108),.res(r36_109),.clk(clk),.wout(w36_109));
	PE pe36_110(.x(x110),.w(w36_109),.acc(r36_109),.res(r36_110),.clk(clk),.wout(w36_110));
	PE pe36_111(.x(x111),.w(w36_110),.acc(r36_110),.res(r36_111),.clk(clk),.wout(w36_111));
	PE pe36_112(.x(x112),.w(w36_111),.acc(r36_111),.res(r36_112),.clk(clk),.wout(w36_112));
	PE pe36_113(.x(x113),.w(w36_112),.acc(r36_112),.res(r36_113),.clk(clk),.wout(w36_113));
	PE pe36_114(.x(x114),.w(w36_113),.acc(r36_113),.res(r36_114),.clk(clk),.wout(w36_114));
	PE pe36_115(.x(x115),.w(w36_114),.acc(r36_114),.res(r36_115),.clk(clk),.wout(w36_115));
	PE pe36_116(.x(x116),.w(w36_115),.acc(r36_115),.res(r36_116),.clk(clk),.wout(w36_116));
	PE pe36_117(.x(x117),.w(w36_116),.acc(r36_116),.res(r36_117),.clk(clk),.wout(w36_117));
	PE pe36_118(.x(x118),.w(w36_117),.acc(r36_117),.res(r36_118),.clk(clk),.wout(w36_118));
	PE pe36_119(.x(x119),.w(w36_118),.acc(r36_118),.res(r36_119),.clk(clk),.wout(w36_119));
	PE pe36_120(.x(x120),.w(w36_119),.acc(r36_119),.res(r36_120),.clk(clk),.wout(w36_120));
	PE pe36_121(.x(x121),.w(w36_120),.acc(r36_120),.res(r36_121),.clk(clk),.wout(w36_121));
	PE pe36_122(.x(x122),.w(w36_121),.acc(r36_121),.res(r36_122),.clk(clk),.wout(w36_122));
	PE pe36_123(.x(x123),.w(w36_122),.acc(r36_122),.res(r36_123),.clk(clk),.wout(w36_123));
	PE pe36_124(.x(x124),.w(w36_123),.acc(r36_123),.res(r36_124),.clk(clk),.wout(w36_124));
	PE pe36_125(.x(x125),.w(w36_124),.acc(r36_124),.res(r36_125),.clk(clk),.wout(w36_125));
	PE pe36_126(.x(x126),.w(w36_125),.acc(r36_125),.res(r36_126),.clk(clk),.wout(w36_126));
	PE pe36_127(.x(x127),.w(w36_126),.acc(r36_126),.res(result36),.clk(clk),.wout(weight36));

	PE pe37_0(.x(x0),.w(w37),.acc(32'h0),.res(r37_0),.clk(clk),.wout(w37_0));
	PE pe37_1(.x(x1),.w(w37_0),.acc(r37_0),.res(r37_1),.clk(clk),.wout(w37_1));
	PE pe37_2(.x(x2),.w(w37_1),.acc(r37_1),.res(r37_2),.clk(clk),.wout(w37_2));
	PE pe37_3(.x(x3),.w(w37_2),.acc(r37_2),.res(r37_3),.clk(clk),.wout(w37_3));
	PE pe37_4(.x(x4),.w(w37_3),.acc(r37_3),.res(r37_4),.clk(clk),.wout(w37_4));
	PE pe37_5(.x(x5),.w(w37_4),.acc(r37_4),.res(r37_5),.clk(clk),.wout(w37_5));
	PE pe37_6(.x(x6),.w(w37_5),.acc(r37_5),.res(r37_6),.clk(clk),.wout(w37_6));
	PE pe37_7(.x(x7),.w(w37_6),.acc(r37_6),.res(r37_7),.clk(clk),.wout(w37_7));
	PE pe37_8(.x(x8),.w(w37_7),.acc(r37_7),.res(r37_8),.clk(clk),.wout(w37_8));
	PE pe37_9(.x(x9),.w(w37_8),.acc(r37_8),.res(r37_9),.clk(clk),.wout(w37_9));
	PE pe37_10(.x(x10),.w(w37_9),.acc(r37_9),.res(r37_10),.clk(clk),.wout(w37_10));
	PE pe37_11(.x(x11),.w(w37_10),.acc(r37_10),.res(r37_11),.clk(clk),.wout(w37_11));
	PE pe37_12(.x(x12),.w(w37_11),.acc(r37_11),.res(r37_12),.clk(clk),.wout(w37_12));
	PE pe37_13(.x(x13),.w(w37_12),.acc(r37_12),.res(r37_13),.clk(clk),.wout(w37_13));
	PE pe37_14(.x(x14),.w(w37_13),.acc(r37_13),.res(r37_14),.clk(clk),.wout(w37_14));
	PE pe37_15(.x(x15),.w(w37_14),.acc(r37_14),.res(r37_15),.clk(clk),.wout(w37_15));
	PE pe37_16(.x(x16),.w(w37_15),.acc(r37_15),.res(r37_16),.clk(clk),.wout(w37_16));
	PE pe37_17(.x(x17),.w(w37_16),.acc(r37_16),.res(r37_17),.clk(clk),.wout(w37_17));
	PE pe37_18(.x(x18),.w(w37_17),.acc(r37_17),.res(r37_18),.clk(clk),.wout(w37_18));
	PE pe37_19(.x(x19),.w(w37_18),.acc(r37_18),.res(r37_19),.clk(clk),.wout(w37_19));
	PE pe37_20(.x(x20),.w(w37_19),.acc(r37_19),.res(r37_20),.clk(clk),.wout(w37_20));
	PE pe37_21(.x(x21),.w(w37_20),.acc(r37_20),.res(r37_21),.clk(clk),.wout(w37_21));
	PE pe37_22(.x(x22),.w(w37_21),.acc(r37_21),.res(r37_22),.clk(clk),.wout(w37_22));
	PE pe37_23(.x(x23),.w(w37_22),.acc(r37_22),.res(r37_23),.clk(clk),.wout(w37_23));
	PE pe37_24(.x(x24),.w(w37_23),.acc(r37_23),.res(r37_24),.clk(clk),.wout(w37_24));
	PE pe37_25(.x(x25),.w(w37_24),.acc(r37_24),.res(r37_25),.clk(clk),.wout(w37_25));
	PE pe37_26(.x(x26),.w(w37_25),.acc(r37_25),.res(r37_26),.clk(clk),.wout(w37_26));
	PE pe37_27(.x(x27),.w(w37_26),.acc(r37_26),.res(r37_27),.clk(clk),.wout(w37_27));
	PE pe37_28(.x(x28),.w(w37_27),.acc(r37_27),.res(r37_28),.clk(clk),.wout(w37_28));
	PE pe37_29(.x(x29),.w(w37_28),.acc(r37_28),.res(r37_29),.clk(clk),.wout(w37_29));
	PE pe37_30(.x(x30),.w(w37_29),.acc(r37_29),.res(r37_30),.clk(clk),.wout(w37_30));
	PE pe37_31(.x(x31),.w(w37_30),.acc(r37_30),.res(r37_31),.clk(clk),.wout(w37_31));
	PE pe37_32(.x(x32),.w(w37_31),.acc(r37_31),.res(r37_32),.clk(clk),.wout(w37_32));
	PE pe37_33(.x(x33),.w(w37_32),.acc(r37_32),.res(r37_33),.clk(clk),.wout(w37_33));
	PE pe37_34(.x(x34),.w(w37_33),.acc(r37_33),.res(r37_34),.clk(clk),.wout(w37_34));
	PE pe37_35(.x(x35),.w(w37_34),.acc(r37_34),.res(r37_35),.clk(clk),.wout(w37_35));
	PE pe37_36(.x(x36),.w(w37_35),.acc(r37_35),.res(r37_36),.clk(clk),.wout(w37_36));
	PE pe37_37(.x(x37),.w(w37_36),.acc(r37_36),.res(r37_37),.clk(clk),.wout(w37_37));
	PE pe37_38(.x(x38),.w(w37_37),.acc(r37_37),.res(r37_38),.clk(clk),.wout(w37_38));
	PE pe37_39(.x(x39),.w(w37_38),.acc(r37_38),.res(r37_39),.clk(clk),.wout(w37_39));
	PE pe37_40(.x(x40),.w(w37_39),.acc(r37_39),.res(r37_40),.clk(clk),.wout(w37_40));
	PE pe37_41(.x(x41),.w(w37_40),.acc(r37_40),.res(r37_41),.clk(clk),.wout(w37_41));
	PE pe37_42(.x(x42),.w(w37_41),.acc(r37_41),.res(r37_42),.clk(clk),.wout(w37_42));
	PE pe37_43(.x(x43),.w(w37_42),.acc(r37_42),.res(r37_43),.clk(clk),.wout(w37_43));
	PE pe37_44(.x(x44),.w(w37_43),.acc(r37_43),.res(r37_44),.clk(clk),.wout(w37_44));
	PE pe37_45(.x(x45),.w(w37_44),.acc(r37_44),.res(r37_45),.clk(clk),.wout(w37_45));
	PE pe37_46(.x(x46),.w(w37_45),.acc(r37_45),.res(r37_46),.clk(clk),.wout(w37_46));
	PE pe37_47(.x(x47),.w(w37_46),.acc(r37_46),.res(r37_47),.clk(clk),.wout(w37_47));
	PE pe37_48(.x(x48),.w(w37_47),.acc(r37_47),.res(r37_48),.clk(clk),.wout(w37_48));
	PE pe37_49(.x(x49),.w(w37_48),.acc(r37_48),.res(r37_49),.clk(clk),.wout(w37_49));
	PE pe37_50(.x(x50),.w(w37_49),.acc(r37_49),.res(r37_50),.clk(clk),.wout(w37_50));
	PE pe37_51(.x(x51),.w(w37_50),.acc(r37_50),.res(r37_51),.clk(clk),.wout(w37_51));
	PE pe37_52(.x(x52),.w(w37_51),.acc(r37_51),.res(r37_52),.clk(clk),.wout(w37_52));
	PE pe37_53(.x(x53),.w(w37_52),.acc(r37_52),.res(r37_53),.clk(clk),.wout(w37_53));
	PE pe37_54(.x(x54),.w(w37_53),.acc(r37_53),.res(r37_54),.clk(clk),.wout(w37_54));
	PE pe37_55(.x(x55),.w(w37_54),.acc(r37_54),.res(r37_55),.clk(clk),.wout(w37_55));
	PE pe37_56(.x(x56),.w(w37_55),.acc(r37_55),.res(r37_56),.clk(clk),.wout(w37_56));
	PE pe37_57(.x(x57),.w(w37_56),.acc(r37_56),.res(r37_57),.clk(clk),.wout(w37_57));
	PE pe37_58(.x(x58),.w(w37_57),.acc(r37_57),.res(r37_58),.clk(clk),.wout(w37_58));
	PE pe37_59(.x(x59),.w(w37_58),.acc(r37_58),.res(r37_59),.clk(clk),.wout(w37_59));
	PE pe37_60(.x(x60),.w(w37_59),.acc(r37_59),.res(r37_60),.clk(clk),.wout(w37_60));
	PE pe37_61(.x(x61),.w(w37_60),.acc(r37_60),.res(r37_61),.clk(clk),.wout(w37_61));
	PE pe37_62(.x(x62),.w(w37_61),.acc(r37_61),.res(r37_62),.clk(clk),.wout(w37_62));
	PE pe37_63(.x(x63),.w(w37_62),.acc(r37_62),.res(r37_63),.clk(clk),.wout(w37_63));
	PE pe37_64(.x(x64),.w(w37_63),.acc(r37_63),.res(r37_64),.clk(clk),.wout(w37_64));
	PE pe37_65(.x(x65),.w(w37_64),.acc(r37_64),.res(r37_65),.clk(clk),.wout(w37_65));
	PE pe37_66(.x(x66),.w(w37_65),.acc(r37_65),.res(r37_66),.clk(clk),.wout(w37_66));
	PE pe37_67(.x(x67),.w(w37_66),.acc(r37_66),.res(r37_67),.clk(clk),.wout(w37_67));
	PE pe37_68(.x(x68),.w(w37_67),.acc(r37_67),.res(r37_68),.clk(clk),.wout(w37_68));
	PE pe37_69(.x(x69),.w(w37_68),.acc(r37_68),.res(r37_69),.clk(clk),.wout(w37_69));
	PE pe37_70(.x(x70),.w(w37_69),.acc(r37_69),.res(r37_70),.clk(clk),.wout(w37_70));
	PE pe37_71(.x(x71),.w(w37_70),.acc(r37_70),.res(r37_71),.clk(clk),.wout(w37_71));
	PE pe37_72(.x(x72),.w(w37_71),.acc(r37_71),.res(r37_72),.clk(clk),.wout(w37_72));
	PE pe37_73(.x(x73),.w(w37_72),.acc(r37_72),.res(r37_73),.clk(clk),.wout(w37_73));
	PE pe37_74(.x(x74),.w(w37_73),.acc(r37_73),.res(r37_74),.clk(clk),.wout(w37_74));
	PE pe37_75(.x(x75),.w(w37_74),.acc(r37_74),.res(r37_75),.clk(clk),.wout(w37_75));
	PE pe37_76(.x(x76),.w(w37_75),.acc(r37_75),.res(r37_76),.clk(clk),.wout(w37_76));
	PE pe37_77(.x(x77),.w(w37_76),.acc(r37_76),.res(r37_77),.clk(clk),.wout(w37_77));
	PE pe37_78(.x(x78),.w(w37_77),.acc(r37_77),.res(r37_78),.clk(clk),.wout(w37_78));
	PE pe37_79(.x(x79),.w(w37_78),.acc(r37_78),.res(r37_79),.clk(clk),.wout(w37_79));
	PE pe37_80(.x(x80),.w(w37_79),.acc(r37_79),.res(r37_80),.clk(clk),.wout(w37_80));
	PE pe37_81(.x(x81),.w(w37_80),.acc(r37_80),.res(r37_81),.clk(clk),.wout(w37_81));
	PE pe37_82(.x(x82),.w(w37_81),.acc(r37_81),.res(r37_82),.clk(clk),.wout(w37_82));
	PE pe37_83(.x(x83),.w(w37_82),.acc(r37_82),.res(r37_83),.clk(clk),.wout(w37_83));
	PE pe37_84(.x(x84),.w(w37_83),.acc(r37_83),.res(r37_84),.clk(clk),.wout(w37_84));
	PE pe37_85(.x(x85),.w(w37_84),.acc(r37_84),.res(r37_85),.clk(clk),.wout(w37_85));
	PE pe37_86(.x(x86),.w(w37_85),.acc(r37_85),.res(r37_86),.clk(clk),.wout(w37_86));
	PE pe37_87(.x(x87),.w(w37_86),.acc(r37_86),.res(r37_87),.clk(clk),.wout(w37_87));
	PE pe37_88(.x(x88),.w(w37_87),.acc(r37_87),.res(r37_88),.clk(clk),.wout(w37_88));
	PE pe37_89(.x(x89),.w(w37_88),.acc(r37_88),.res(r37_89),.clk(clk),.wout(w37_89));
	PE pe37_90(.x(x90),.w(w37_89),.acc(r37_89),.res(r37_90),.clk(clk),.wout(w37_90));
	PE pe37_91(.x(x91),.w(w37_90),.acc(r37_90),.res(r37_91),.clk(clk),.wout(w37_91));
	PE pe37_92(.x(x92),.w(w37_91),.acc(r37_91),.res(r37_92),.clk(clk),.wout(w37_92));
	PE pe37_93(.x(x93),.w(w37_92),.acc(r37_92),.res(r37_93),.clk(clk),.wout(w37_93));
	PE pe37_94(.x(x94),.w(w37_93),.acc(r37_93),.res(r37_94),.clk(clk),.wout(w37_94));
	PE pe37_95(.x(x95),.w(w37_94),.acc(r37_94),.res(r37_95),.clk(clk),.wout(w37_95));
	PE pe37_96(.x(x96),.w(w37_95),.acc(r37_95),.res(r37_96),.clk(clk),.wout(w37_96));
	PE pe37_97(.x(x97),.w(w37_96),.acc(r37_96),.res(r37_97),.clk(clk),.wout(w37_97));
	PE pe37_98(.x(x98),.w(w37_97),.acc(r37_97),.res(r37_98),.clk(clk),.wout(w37_98));
	PE pe37_99(.x(x99),.w(w37_98),.acc(r37_98),.res(r37_99),.clk(clk),.wout(w37_99));
	PE pe37_100(.x(x100),.w(w37_99),.acc(r37_99),.res(r37_100),.clk(clk),.wout(w37_100));
	PE pe37_101(.x(x101),.w(w37_100),.acc(r37_100),.res(r37_101),.clk(clk),.wout(w37_101));
	PE pe37_102(.x(x102),.w(w37_101),.acc(r37_101),.res(r37_102),.clk(clk),.wout(w37_102));
	PE pe37_103(.x(x103),.w(w37_102),.acc(r37_102),.res(r37_103),.clk(clk),.wout(w37_103));
	PE pe37_104(.x(x104),.w(w37_103),.acc(r37_103),.res(r37_104),.clk(clk),.wout(w37_104));
	PE pe37_105(.x(x105),.w(w37_104),.acc(r37_104),.res(r37_105),.clk(clk),.wout(w37_105));
	PE pe37_106(.x(x106),.w(w37_105),.acc(r37_105),.res(r37_106),.clk(clk),.wout(w37_106));
	PE pe37_107(.x(x107),.w(w37_106),.acc(r37_106),.res(r37_107),.clk(clk),.wout(w37_107));
	PE pe37_108(.x(x108),.w(w37_107),.acc(r37_107),.res(r37_108),.clk(clk),.wout(w37_108));
	PE pe37_109(.x(x109),.w(w37_108),.acc(r37_108),.res(r37_109),.clk(clk),.wout(w37_109));
	PE pe37_110(.x(x110),.w(w37_109),.acc(r37_109),.res(r37_110),.clk(clk),.wout(w37_110));
	PE pe37_111(.x(x111),.w(w37_110),.acc(r37_110),.res(r37_111),.clk(clk),.wout(w37_111));
	PE pe37_112(.x(x112),.w(w37_111),.acc(r37_111),.res(r37_112),.clk(clk),.wout(w37_112));
	PE pe37_113(.x(x113),.w(w37_112),.acc(r37_112),.res(r37_113),.clk(clk),.wout(w37_113));
	PE pe37_114(.x(x114),.w(w37_113),.acc(r37_113),.res(r37_114),.clk(clk),.wout(w37_114));
	PE pe37_115(.x(x115),.w(w37_114),.acc(r37_114),.res(r37_115),.clk(clk),.wout(w37_115));
	PE pe37_116(.x(x116),.w(w37_115),.acc(r37_115),.res(r37_116),.clk(clk),.wout(w37_116));
	PE pe37_117(.x(x117),.w(w37_116),.acc(r37_116),.res(r37_117),.clk(clk),.wout(w37_117));
	PE pe37_118(.x(x118),.w(w37_117),.acc(r37_117),.res(r37_118),.clk(clk),.wout(w37_118));
	PE pe37_119(.x(x119),.w(w37_118),.acc(r37_118),.res(r37_119),.clk(clk),.wout(w37_119));
	PE pe37_120(.x(x120),.w(w37_119),.acc(r37_119),.res(r37_120),.clk(clk),.wout(w37_120));
	PE pe37_121(.x(x121),.w(w37_120),.acc(r37_120),.res(r37_121),.clk(clk),.wout(w37_121));
	PE pe37_122(.x(x122),.w(w37_121),.acc(r37_121),.res(r37_122),.clk(clk),.wout(w37_122));
	PE pe37_123(.x(x123),.w(w37_122),.acc(r37_122),.res(r37_123),.clk(clk),.wout(w37_123));
	PE pe37_124(.x(x124),.w(w37_123),.acc(r37_123),.res(r37_124),.clk(clk),.wout(w37_124));
	PE pe37_125(.x(x125),.w(w37_124),.acc(r37_124),.res(r37_125),.clk(clk),.wout(w37_125));
	PE pe37_126(.x(x126),.w(w37_125),.acc(r37_125),.res(r37_126),.clk(clk),.wout(w37_126));
	PE pe37_127(.x(x127),.w(w37_126),.acc(r37_126),.res(result37),.clk(clk),.wout(weight37));

	PE pe38_0(.x(x0),.w(w38),.acc(32'h0),.res(r38_0),.clk(clk),.wout(w38_0));
	PE pe38_1(.x(x1),.w(w38_0),.acc(r38_0),.res(r38_1),.clk(clk),.wout(w38_1));
	PE pe38_2(.x(x2),.w(w38_1),.acc(r38_1),.res(r38_2),.clk(clk),.wout(w38_2));
	PE pe38_3(.x(x3),.w(w38_2),.acc(r38_2),.res(r38_3),.clk(clk),.wout(w38_3));
	PE pe38_4(.x(x4),.w(w38_3),.acc(r38_3),.res(r38_4),.clk(clk),.wout(w38_4));
	PE pe38_5(.x(x5),.w(w38_4),.acc(r38_4),.res(r38_5),.clk(clk),.wout(w38_5));
	PE pe38_6(.x(x6),.w(w38_5),.acc(r38_5),.res(r38_6),.clk(clk),.wout(w38_6));
	PE pe38_7(.x(x7),.w(w38_6),.acc(r38_6),.res(r38_7),.clk(clk),.wout(w38_7));
	PE pe38_8(.x(x8),.w(w38_7),.acc(r38_7),.res(r38_8),.clk(clk),.wout(w38_8));
	PE pe38_9(.x(x9),.w(w38_8),.acc(r38_8),.res(r38_9),.clk(clk),.wout(w38_9));
	PE pe38_10(.x(x10),.w(w38_9),.acc(r38_9),.res(r38_10),.clk(clk),.wout(w38_10));
	PE pe38_11(.x(x11),.w(w38_10),.acc(r38_10),.res(r38_11),.clk(clk),.wout(w38_11));
	PE pe38_12(.x(x12),.w(w38_11),.acc(r38_11),.res(r38_12),.clk(clk),.wout(w38_12));
	PE pe38_13(.x(x13),.w(w38_12),.acc(r38_12),.res(r38_13),.clk(clk),.wout(w38_13));
	PE pe38_14(.x(x14),.w(w38_13),.acc(r38_13),.res(r38_14),.clk(clk),.wout(w38_14));
	PE pe38_15(.x(x15),.w(w38_14),.acc(r38_14),.res(r38_15),.clk(clk),.wout(w38_15));
	PE pe38_16(.x(x16),.w(w38_15),.acc(r38_15),.res(r38_16),.clk(clk),.wout(w38_16));
	PE pe38_17(.x(x17),.w(w38_16),.acc(r38_16),.res(r38_17),.clk(clk),.wout(w38_17));
	PE pe38_18(.x(x18),.w(w38_17),.acc(r38_17),.res(r38_18),.clk(clk),.wout(w38_18));
	PE pe38_19(.x(x19),.w(w38_18),.acc(r38_18),.res(r38_19),.clk(clk),.wout(w38_19));
	PE pe38_20(.x(x20),.w(w38_19),.acc(r38_19),.res(r38_20),.clk(clk),.wout(w38_20));
	PE pe38_21(.x(x21),.w(w38_20),.acc(r38_20),.res(r38_21),.clk(clk),.wout(w38_21));
	PE pe38_22(.x(x22),.w(w38_21),.acc(r38_21),.res(r38_22),.clk(clk),.wout(w38_22));
	PE pe38_23(.x(x23),.w(w38_22),.acc(r38_22),.res(r38_23),.clk(clk),.wout(w38_23));
	PE pe38_24(.x(x24),.w(w38_23),.acc(r38_23),.res(r38_24),.clk(clk),.wout(w38_24));
	PE pe38_25(.x(x25),.w(w38_24),.acc(r38_24),.res(r38_25),.clk(clk),.wout(w38_25));
	PE pe38_26(.x(x26),.w(w38_25),.acc(r38_25),.res(r38_26),.clk(clk),.wout(w38_26));
	PE pe38_27(.x(x27),.w(w38_26),.acc(r38_26),.res(r38_27),.clk(clk),.wout(w38_27));
	PE pe38_28(.x(x28),.w(w38_27),.acc(r38_27),.res(r38_28),.clk(clk),.wout(w38_28));
	PE pe38_29(.x(x29),.w(w38_28),.acc(r38_28),.res(r38_29),.clk(clk),.wout(w38_29));
	PE pe38_30(.x(x30),.w(w38_29),.acc(r38_29),.res(r38_30),.clk(clk),.wout(w38_30));
	PE pe38_31(.x(x31),.w(w38_30),.acc(r38_30),.res(r38_31),.clk(clk),.wout(w38_31));
	PE pe38_32(.x(x32),.w(w38_31),.acc(r38_31),.res(r38_32),.clk(clk),.wout(w38_32));
	PE pe38_33(.x(x33),.w(w38_32),.acc(r38_32),.res(r38_33),.clk(clk),.wout(w38_33));
	PE pe38_34(.x(x34),.w(w38_33),.acc(r38_33),.res(r38_34),.clk(clk),.wout(w38_34));
	PE pe38_35(.x(x35),.w(w38_34),.acc(r38_34),.res(r38_35),.clk(clk),.wout(w38_35));
	PE pe38_36(.x(x36),.w(w38_35),.acc(r38_35),.res(r38_36),.clk(clk),.wout(w38_36));
	PE pe38_37(.x(x37),.w(w38_36),.acc(r38_36),.res(r38_37),.clk(clk),.wout(w38_37));
	PE pe38_38(.x(x38),.w(w38_37),.acc(r38_37),.res(r38_38),.clk(clk),.wout(w38_38));
	PE pe38_39(.x(x39),.w(w38_38),.acc(r38_38),.res(r38_39),.clk(clk),.wout(w38_39));
	PE pe38_40(.x(x40),.w(w38_39),.acc(r38_39),.res(r38_40),.clk(clk),.wout(w38_40));
	PE pe38_41(.x(x41),.w(w38_40),.acc(r38_40),.res(r38_41),.clk(clk),.wout(w38_41));
	PE pe38_42(.x(x42),.w(w38_41),.acc(r38_41),.res(r38_42),.clk(clk),.wout(w38_42));
	PE pe38_43(.x(x43),.w(w38_42),.acc(r38_42),.res(r38_43),.clk(clk),.wout(w38_43));
	PE pe38_44(.x(x44),.w(w38_43),.acc(r38_43),.res(r38_44),.clk(clk),.wout(w38_44));
	PE pe38_45(.x(x45),.w(w38_44),.acc(r38_44),.res(r38_45),.clk(clk),.wout(w38_45));
	PE pe38_46(.x(x46),.w(w38_45),.acc(r38_45),.res(r38_46),.clk(clk),.wout(w38_46));
	PE pe38_47(.x(x47),.w(w38_46),.acc(r38_46),.res(r38_47),.clk(clk),.wout(w38_47));
	PE pe38_48(.x(x48),.w(w38_47),.acc(r38_47),.res(r38_48),.clk(clk),.wout(w38_48));
	PE pe38_49(.x(x49),.w(w38_48),.acc(r38_48),.res(r38_49),.clk(clk),.wout(w38_49));
	PE pe38_50(.x(x50),.w(w38_49),.acc(r38_49),.res(r38_50),.clk(clk),.wout(w38_50));
	PE pe38_51(.x(x51),.w(w38_50),.acc(r38_50),.res(r38_51),.clk(clk),.wout(w38_51));
	PE pe38_52(.x(x52),.w(w38_51),.acc(r38_51),.res(r38_52),.clk(clk),.wout(w38_52));
	PE pe38_53(.x(x53),.w(w38_52),.acc(r38_52),.res(r38_53),.clk(clk),.wout(w38_53));
	PE pe38_54(.x(x54),.w(w38_53),.acc(r38_53),.res(r38_54),.clk(clk),.wout(w38_54));
	PE pe38_55(.x(x55),.w(w38_54),.acc(r38_54),.res(r38_55),.clk(clk),.wout(w38_55));
	PE pe38_56(.x(x56),.w(w38_55),.acc(r38_55),.res(r38_56),.clk(clk),.wout(w38_56));
	PE pe38_57(.x(x57),.w(w38_56),.acc(r38_56),.res(r38_57),.clk(clk),.wout(w38_57));
	PE pe38_58(.x(x58),.w(w38_57),.acc(r38_57),.res(r38_58),.clk(clk),.wout(w38_58));
	PE pe38_59(.x(x59),.w(w38_58),.acc(r38_58),.res(r38_59),.clk(clk),.wout(w38_59));
	PE pe38_60(.x(x60),.w(w38_59),.acc(r38_59),.res(r38_60),.clk(clk),.wout(w38_60));
	PE pe38_61(.x(x61),.w(w38_60),.acc(r38_60),.res(r38_61),.clk(clk),.wout(w38_61));
	PE pe38_62(.x(x62),.w(w38_61),.acc(r38_61),.res(r38_62),.clk(clk),.wout(w38_62));
	PE pe38_63(.x(x63),.w(w38_62),.acc(r38_62),.res(r38_63),.clk(clk),.wout(w38_63));
	PE pe38_64(.x(x64),.w(w38_63),.acc(r38_63),.res(r38_64),.clk(clk),.wout(w38_64));
	PE pe38_65(.x(x65),.w(w38_64),.acc(r38_64),.res(r38_65),.clk(clk),.wout(w38_65));
	PE pe38_66(.x(x66),.w(w38_65),.acc(r38_65),.res(r38_66),.clk(clk),.wout(w38_66));
	PE pe38_67(.x(x67),.w(w38_66),.acc(r38_66),.res(r38_67),.clk(clk),.wout(w38_67));
	PE pe38_68(.x(x68),.w(w38_67),.acc(r38_67),.res(r38_68),.clk(clk),.wout(w38_68));
	PE pe38_69(.x(x69),.w(w38_68),.acc(r38_68),.res(r38_69),.clk(clk),.wout(w38_69));
	PE pe38_70(.x(x70),.w(w38_69),.acc(r38_69),.res(r38_70),.clk(clk),.wout(w38_70));
	PE pe38_71(.x(x71),.w(w38_70),.acc(r38_70),.res(r38_71),.clk(clk),.wout(w38_71));
	PE pe38_72(.x(x72),.w(w38_71),.acc(r38_71),.res(r38_72),.clk(clk),.wout(w38_72));
	PE pe38_73(.x(x73),.w(w38_72),.acc(r38_72),.res(r38_73),.clk(clk),.wout(w38_73));
	PE pe38_74(.x(x74),.w(w38_73),.acc(r38_73),.res(r38_74),.clk(clk),.wout(w38_74));
	PE pe38_75(.x(x75),.w(w38_74),.acc(r38_74),.res(r38_75),.clk(clk),.wout(w38_75));
	PE pe38_76(.x(x76),.w(w38_75),.acc(r38_75),.res(r38_76),.clk(clk),.wout(w38_76));
	PE pe38_77(.x(x77),.w(w38_76),.acc(r38_76),.res(r38_77),.clk(clk),.wout(w38_77));
	PE pe38_78(.x(x78),.w(w38_77),.acc(r38_77),.res(r38_78),.clk(clk),.wout(w38_78));
	PE pe38_79(.x(x79),.w(w38_78),.acc(r38_78),.res(r38_79),.clk(clk),.wout(w38_79));
	PE pe38_80(.x(x80),.w(w38_79),.acc(r38_79),.res(r38_80),.clk(clk),.wout(w38_80));
	PE pe38_81(.x(x81),.w(w38_80),.acc(r38_80),.res(r38_81),.clk(clk),.wout(w38_81));
	PE pe38_82(.x(x82),.w(w38_81),.acc(r38_81),.res(r38_82),.clk(clk),.wout(w38_82));
	PE pe38_83(.x(x83),.w(w38_82),.acc(r38_82),.res(r38_83),.clk(clk),.wout(w38_83));
	PE pe38_84(.x(x84),.w(w38_83),.acc(r38_83),.res(r38_84),.clk(clk),.wout(w38_84));
	PE pe38_85(.x(x85),.w(w38_84),.acc(r38_84),.res(r38_85),.clk(clk),.wout(w38_85));
	PE pe38_86(.x(x86),.w(w38_85),.acc(r38_85),.res(r38_86),.clk(clk),.wout(w38_86));
	PE pe38_87(.x(x87),.w(w38_86),.acc(r38_86),.res(r38_87),.clk(clk),.wout(w38_87));
	PE pe38_88(.x(x88),.w(w38_87),.acc(r38_87),.res(r38_88),.clk(clk),.wout(w38_88));
	PE pe38_89(.x(x89),.w(w38_88),.acc(r38_88),.res(r38_89),.clk(clk),.wout(w38_89));
	PE pe38_90(.x(x90),.w(w38_89),.acc(r38_89),.res(r38_90),.clk(clk),.wout(w38_90));
	PE pe38_91(.x(x91),.w(w38_90),.acc(r38_90),.res(r38_91),.clk(clk),.wout(w38_91));
	PE pe38_92(.x(x92),.w(w38_91),.acc(r38_91),.res(r38_92),.clk(clk),.wout(w38_92));
	PE pe38_93(.x(x93),.w(w38_92),.acc(r38_92),.res(r38_93),.clk(clk),.wout(w38_93));
	PE pe38_94(.x(x94),.w(w38_93),.acc(r38_93),.res(r38_94),.clk(clk),.wout(w38_94));
	PE pe38_95(.x(x95),.w(w38_94),.acc(r38_94),.res(r38_95),.clk(clk),.wout(w38_95));
	PE pe38_96(.x(x96),.w(w38_95),.acc(r38_95),.res(r38_96),.clk(clk),.wout(w38_96));
	PE pe38_97(.x(x97),.w(w38_96),.acc(r38_96),.res(r38_97),.clk(clk),.wout(w38_97));
	PE pe38_98(.x(x98),.w(w38_97),.acc(r38_97),.res(r38_98),.clk(clk),.wout(w38_98));
	PE pe38_99(.x(x99),.w(w38_98),.acc(r38_98),.res(r38_99),.clk(clk),.wout(w38_99));
	PE pe38_100(.x(x100),.w(w38_99),.acc(r38_99),.res(r38_100),.clk(clk),.wout(w38_100));
	PE pe38_101(.x(x101),.w(w38_100),.acc(r38_100),.res(r38_101),.clk(clk),.wout(w38_101));
	PE pe38_102(.x(x102),.w(w38_101),.acc(r38_101),.res(r38_102),.clk(clk),.wout(w38_102));
	PE pe38_103(.x(x103),.w(w38_102),.acc(r38_102),.res(r38_103),.clk(clk),.wout(w38_103));
	PE pe38_104(.x(x104),.w(w38_103),.acc(r38_103),.res(r38_104),.clk(clk),.wout(w38_104));
	PE pe38_105(.x(x105),.w(w38_104),.acc(r38_104),.res(r38_105),.clk(clk),.wout(w38_105));
	PE pe38_106(.x(x106),.w(w38_105),.acc(r38_105),.res(r38_106),.clk(clk),.wout(w38_106));
	PE pe38_107(.x(x107),.w(w38_106),.acc(r38_106),.res(r38_107),.clk(clk),.wout(w38_107));
	PE pe38_108(.x(x108),.w(w38_107),.acc(r38_107),.res(r38_108),.clk(clk),.wout(w38_108));
	PE pe38_109(.x(x109),.w(w38_108),.acc(r38_108),.res(r38_109),.clk(clk),.wout(w38_109));
	PE pe38_110(.x(x110),.w(w38_109),.acc(r38_109),.res(r38_110),.clk(clk),.wout(w38_110));
	PE pe38_111(.x(x111),.w(w38_110),.acc(r38_110),.res(r38_111),.clk(clk),.wout(w38_111));
	PE pe38_112(.x(x112),.w(w38_111),.acc(r38_111),.res(r38_112),.clk(clk),.wout(w38_112));
	PE pe38_113(.x(x113),.w(w38_112),.acc(r38_112),.res(r38_113),.clk(clk),.wout(w38_113));
	PE pe38_114(.x(x114),.w(w38_113),.acc(r38_113),.res(r38_114),.clk(clk),.wout(w38_114));
	PE pe38_115(.x(x115),.w(w38_114),.acc(r38_114),.res(r38_115),.clk(clk),.wout(w38_115));
	PE pe38_116(.x(x116),.w(w38_115),.acc(r38_115),.res(r38_116),.clk(clk),.wout(w38_116));
	PE pe38_117(.x(x117),.w(w38_116),.acc(r38_116),.res(r38_117),.clk(clk),.wout(w38_117));
	PE pe38_118(.x(x118),.w(w38_117),.acc(r38_117),.res(r38_118),.clk(clk),.wout(w38_118));
	PE pe38_119(.x(x119),.w(w38_118),.acc(r38_118),.res(r38_119),.clk(clk),.wout(w38_119));
	PE pe38_120(.x(x120),.w(w38_119),.acc(r38_119),.res(r38_120),.clk(clk),.wout(w38_120));
	PE pe38_121(.x(x121),.w(w38_120),.acc(r38_120),.res(r38_121),.clk(clk),.wout(w38_121));
	PE pe38_122(.x(x122),.w(w38_121),.acc(r38_121),.res(r38_122),.clk(clk),.wout(w38_122));
	PE pe38_123(.x(x123),.w(w38_122),.acc(r38_122),.res(r38_123),.clk(clk),.wout(w38_123));
	PE pe38_124(.x(x124),.w(w38_123),.acc(r38_123),.res(r38_124),.clk(clk),.wout(w38_124));
	PE pe38_125(.x(x125),.w(w38_124),.acc(r38_124),.res(r38_125),.clk(clk),.wout(w38_125));
	PE pe38_126(.x(x126),.w(w38_125),.acc(r38_125),.res(r38_126),.clk(clk),.wout(w38_126));
	PE pe38_127(.x(x127),.w(w38_126),.acc(r38_126),.res(result38),.clk(clk),.wout(weight38));

	PE pe39_0(.x(x0),.w(w39),.acc(32'h0),.res(r39_0),.clk(clk),.wout(w39_0));
	PE pe39_1(.x(x1),.w(w39_0),.acc(r39_0),.res(r39_1),.clk(clk),.wout(w39_1));
	PE pe39_2(.x(x2),.w(w39_1),.acc(r39_1),.res(r39_2),.clk(clk),.wout(w39_2));
	PE pe39_3(.x(x3),.w(w39_2),.acc(r39_2),.res(r39_3),.clk(clk),.wout(w39_3));
	PE pe39_4(.x(x4),.w(w39_3),.acc(r39_3),.res(r39_4),.clk(clk),.wout(w39_4));
	PE pe39_5(.x(x5),.w(w39_4),.acc(r39_4),.res(r39_5),.clk(clk),.wout(w39_5));
	PE pe39_6(.x(x6),.w(w39_5),.acc(r39_5),.res(r39_6),.clk(clk),.wout(w39_6));
	PE pe39_7(.x(x7),.w(w39_6),.acc(r39_6),.res(r39_7),.clk(clk),.wout(w39_7));
	PE pe39_8(.x(x8),.w(w39_7),.acc(r39_7),.res(r39_8),.clk(clk),.wout(w39_8));
	PE pe39_9(.x(x9),.w(w39_8),.acc(r39_8),.res(r39_9),.clk(clk),.wout(w39_9));
	PE pe39_10(.x(x10),.w(w39_9),.acc(r39_9),.res(r39_10),.clk(clk),.wout(w39_10));
	PE pe39_11(.x(x11),.w(w39_10),.acc(r39_10),.res(r39_11),.clk(clk),.wout(w39_11));
	PE pe39_12(.x(x12),.w(w39_11),.acc(r39_11),.res(r39_12),.clk(clk),.wout(w39_12));
	PE pe39_13(.x(x13),.w(w39_12),.acc(r39_12),.res(r39_13),.clk(clk),.wout(w39_13));
	PE pe39_14(.x(x14),.w(w39_13),.acc(r39_13),.res(r39_14),.clk(clk),.wout(w39_14));
	PE pe39_15(.x(x15),.w(w39_14),.acc(r39_14),.res(r39_15),.clk(clk),.wout(w39_15));
	PE pe39_16(.x(x16),.w(w39_15),.acc(r39_15),.res(r39_16),.clk(clk),.wout(w39_16));
	PE pe39_17(.x(x17),.w(w39_16),.acc(r39_16),.res(r39_17),.clk(clk),.wout(w39_17));
	PE pe39_18(.x(x18),.w(w39_17),.acc(r39_17),.res(r39_18),.clk(clk),.wout(w39_18));
	PE pe39_19(.x(x19),.w(w39_18),.acc(r39_18),.res(r39_19),.clk(clk),.wout(w39_19));
	PE pe39_20(.x(x20),.w(w39_19),.acc(r39_19),.res(r39_20),.clk(clk),.wout(w39_20));
	PE pe39_21(.x(x21),.w(w39_20),.acc(r39_20),.res(r39_21),.clk(clk),.wout(w39_21));
	PE pe39_22(.x(x22),.w(w39_21),.acc(r39_21),.res(r39_22),.clk(clk),.wout(w39_22));
	PE pe39_23(.x(x23),.w(w39_22),.acc(r39_22),.res(r39_23),.clk(clk),.wout(w39_23));
	PE pe39_24(.x(x24),.w(w39_23),.acc(r39_23),.res(r39_24),.clk(clk),.wout(w39_24));
	PE pe39_25(.x(x25),.w(w39_24),.acc(r39_24),.res(r39_25),.clk(clk),.wout(w39_25));
	PE pe39_26(.x(x26),.w(w39_25),.acc(r39_25),.res(r39_26),.clk(clk),.wout(w39_26));
	PE pe39_27(.x(x27),.w(w39_26),.acc(r39_26),.res(r39_27),.clk(clk),.wout(w39_27));
	PE pe39_28(.x(x28),.w(w39_27),.acc(r39_27),.res(r39_28),.clk(clk),.wout(w39_28));
	PE pe39_29(.x(x29),.w(w39_28),.acc(r39_28),.res(r39_29),.clk(clk),.wout(w39_29));
	PE pe39_30(.x(x30),.w(w39_29),.acc(r39_29),.res(r39_30),.clk(clk),.wout(w39_30));
	PE pe39_31(.x(x31),.w(w39_30),.acc(r39_30),.res(r39_31),.clk(clk),.wout(w39_31));
	PE pe39_32(.x(x32),.w(w39_31),.acc(r39_31),.res(r39_32),.clk(clk),.wout(w39_32));
	PE pe39_33(.x(x33),.w(w39_32),.acc(r39_32),.res(r39_33),.clk(clk),.wout(w39_33));
	PE pe39_34(.x(x34),.w(w39_33),.acc(r39_33),.res(r39_34),.clk(clk),.wout(w39_34));
	PE pe39_35(.x(x35),.w(w39_34),.acc(r39_34),.res(r39_35),.clk(clk),.wout(w39_35));
	PE pe39_36(.x(x36),.w(w39_35),.acc(r39_35),.res(r39_36),.clk(clk),.wout(w39_36));
	PE pe39_37(.x(x37),.w(w39_36),.acc(r39_36),.res(r39_37),.clk(clk),.wout(w39_37));
	PE pe39_38(.x(x38),.w(w39_37),.acc(r39_37),.res(r39_38),.clk(clk),.wout(w39_38));
	PE pe39_39(.x(x39),.w(w39_38),.acc(r39_38),.res(r39_39),.clk(clk),.wout(w39_39));
	PE pe39_40(.x(x40),.w(w39_39),.acc(r39_39),.res(r39_40),.clk(clk),.wout(w39_40));
	PE pe39_41(.x(x41),.w(w39_40),.acc(r39_40),.res(r39_41),.clk(clk),.wout(w39_41));
	PE pe39_42(.x(x42),.w(w39_41),.acc(r39_41),.res(r39_42),.clk(clk),.wout(w39_42));
	PE pe39_43(.x(x43),.w(w39_42),.acc(r39_42),.res(r39_43),.clk(clk),.wout(w39_43));
	PE pe39_44(.x(x44),.w(w39_43),.acc(r39_43),.res(r39_44),.clk(clk),.wout(w39_44));
	PE pe39_45(.x(x45),.w(w39_44),.acc(r39_44),.res(r39_45),.clk(clk),.wout(w39_45));
	PE pe39_46(.x(x46),.w(w39_45),.acc(r39_45),.res(r39_46),.clk(clk),.wout(w39_46));
	PE pe39_47(.x(x47),.w(w39_46),.acc(r39_46),.res(r39_47),.clk(clk),.wout(w39_47));
	PE pe39_48(.x(x48),.w(w39_47),.acc(r39_47),.res(r39_48),.clk(clk),.wout(w39_48));
	PE pe39_49(.x(x49),.w(w39_48),.acc(r39_48),.res(r39_49),.clk(clk),.wout(w39_49));
	PE pe39_50(.x(x50),.w(w39_49),.acc(r39_49),.res(r39_50),.clk(clk),.wout(w39_50));
	PE pe39_51(.x(x51),.w(w39_50),.acc(r39_50),.res(r39_51),.clk(clk),.wout(w39_51));
	PE pe39_52(.x(x52),.w(w39_51),.acc(r39_51),.res(r39_52),.clk(clk),.wout(w39_52));
	PE pe39_53(.x(x53),.w(w39_52),.acc(r39_52),.res(r39_53),.clk(clk),.wout(w39_53));
	PE pe39_54(.x(x54),.w(w39_53),.acc(r39_53),.res(r39_54),.clk(clk),.wout(w39_54));
	PE pe39_55(.x(x55),.w(w39_54),.acc(r39_54),.res(r39_55),.clk(clk),.wout(w39_55));
	PE pe39_56(.x(x56),.w(w39_55),.acc(r39_55),.res(r39_56),.clk(clk),.wout(w39_56));
	PE pe39_57(.x(x57),.w(w39_56),.acc(r39_56),.res(r39_57),.clk(clk),.wout(w39_57));
	PE pe39_58(.x(x58),.w(w39_57),.acc(r39_57),.res(r39_58),.clk(clk),.wout(w39_58));
	PE pe39_59(.x(x59),.w(w39_58),.acc(r39_58),.res(r39_59),.clk(clk),.wout(w39_59));
	PE pe39_60(.x(x60),.w(w39_59),.acc(r39_59),.res(r39_60),.clk(clk),.wout(w39_60));
	PE pe39_61(.x(x61),.w(w39_60),.acc(r39_60),.res(r39_61),.clk(clk),.wout(w39_61));
	PE pe39_62(.x(x62),.w(w39_61),.acc(r39_61),.res(r39_62),.clk(clk),.wout(w39_62));
	PE pe39_63(.x(x63),.w(w39_62),.acc(r39_62),.res(r39_63),.clk(clk),.wout(w39_63));
	PE pe39_64(.x(x64),.w(w39_63),.acc(r39_63),.res(r39_64),.clk(clk),.wout(w39_64));
	PE pe39_65(.x(x65),.w(w39_64),.acc(r39_64),.res(r39_65),.clk(clk),.wout(w39_65));
	PE pe39_66(.x(x66),.w(w39_65),.acc(r39_65),.res(r39_66),.clk(clk),.wout(w39_66));
	PE pe39_67(.x(x67),.w(w39_66),.acc(r39_66),.res(r39_67),.clk(clk),.wout(w39_67));
	PE pe39_68(.x(x68),.w(w39_67),.acc(r39_67),.res(r39_68),.clk(clk),.wout(w39_68));
	PE pe39_69(.x(x69),.w(w39_68),.acc(r39_68),.res(r39_69),.clk(clk),.wout(w39_69));
	PE pe39_70(.x(x70),.w(w39_69),.acc(r39_69),.res(r39_70),.clk(clk),.wout(w39_70));
	PE pe39_71(.x(x71),.w(w39_70),.acc(r39_70),.res(r39_71),.clk(clk),.wout(w39_71));
	PE pe39_72(.x(x72),.w(w39_71),.acc(r39_71),.res(r39_72),.clk(clk),.wout(w39_72));
	PE pe39_73(.x(x73),.w(w39_72),.acc(r39_72),.res(r39_73),.clk(clk),.wout(w39_73));
	PE pe39_74(.x(x74),.w(w39_73),.acc(r39_73),.res(r39_74),.clk(clk),.wout(w39_74));
	PE pe39_75(.x(x75),.w(w39_74),.acc(r39_74),.res(r39_75),.clk(clk),.wout(w39_75));
	PE pe39_76(.x(x76),.w(w39_75),.acc(r39_75),.res(r39_76),.clk(clk),.wout(w39_76));
	PE pe39_77(.x(x77),.w(w39_76),.acc(r39_76),.res(r39_77),.clk(clk),.wout(w39_77));
	PE pe39_78(.x(x78),.w(w39_77),.acc(r39_77),.res(r39_78),.clk(clk),.wout(w39_78));
	PE pe39_79(.x(x79),.w(w39_78),.acc(r39_78),.res(r39_79),.clk(clk),.wout(w39_79));
	PE pe39_80(.x(x80),.w(w39_79),.acc(r39_79),.res(r39_80),.clk(clk),.wout(w39_80));
	PE pe39_81(.x(x81),.w(w39_80),.acc(r39_80),.res(r39_81),.clk(clk),.wout(w39_81));
	PE pe39_82(.x(x82),.w(w39_81),.acc(r39_81),.res(r39_82),.clk(clk),.wout(w39_82));
	PE pe39_83(.x(x83),.w(w39_82),.acc(r39_82),.res(r39_83),.clk(clk),.wout(w39_83));
	PE pe39_84(.x(x84),.w(w39_83),.acc(r39_83),.res(r39_84),.clk(clk),.wout(w39_84));
	PE pe39_85(.x(x85),.w(w39_84),.acc(r39_84),.res(r39_85),.clk(clk),.wout(w39_85));
	PE pe39_86(.x(x86),.w(w39_85),.acc(r39_85),.res(r39_86),.clk(clk),.wout(w39_86));
	PE pe39_87(.x(x87),.w(w39_86),.acc(r39_86),.res(r39_87),.clk(clk),.wout(w39_87));
	PE pe39_88(.x(x88),.w(w39_87),.acc(r39_87),.res(r39_88),.clk(clk),.wout(w39_88));
	PE pe39_89(.x(x89),.w(w39_88),.acc(r39_88),.res(r39_89),.clk(clk),.wout(w39_89));
	PE pe39_90(.x(x90),.w(w39_89),.acc(r39_89),.res(r39_90),.clk(clk),.wout(w39_90));
	PE pe39_91(.x(x91),.w(w39_90),.acc(r39_90),.res(r39_91),.clk(clk),.wout(w39_91));
	PE pe39_92(.x(x92),.w(w39_91),.acc(r39_91),.res(r39_92),.clk(clk),.wout(w39_92));
	PE pe39_93(.x(x93),.w(w39_92),.acc(r39_92),.res(r39_93),.clk(clk),.wout(w39_93));
	PE pe39_94(.x(x94),.w(w39_93),.acc(r39_93),.res(r39_94),.clk(clk),.wout(w39_94));
	PE pe39_95(.x(x95),.w(w39_94),.acc(r39_94),.res(r39_95),.clk(clk),.wout(w39_95));
	PE pe39_96(.x(x96),.w(w39_95),.acc(r39_95),.res(r39_96),.clk(clk),.wout(w39_96));
	PE pe39_97(.x(x97),.w(w39_96),.acc(r39_96),.res(r39_97),.clk(clk),.wout(w39_97));
	PE pe39_98(.x(x98),.w(w39_97),.acc(r39_97),.res(r39_98),.clk(clk),.wout(w39_98));
	PE pe39_99(.x(x99),.w(w39_98),.acc(r39_98),.res(r39_99),.clk(clk),.wout(w39_99));
	PE pe39_100(.x(x100),.w(w39_99),.acc(r39_99),.res(r39_100),.clk(clk),.wout(w39_100));
	PE pe39_101(.x(x101),.w(w39_100),.acc(r39_100),.res(r39_101),.clk(clk),.wout(w39_101));
	PE pe39_102(.x(x102),.w(w39_101),.acc(r39_101),.res(r39_102),.clk(clk),.wout(w39_102));
	PE pe39_103(.x(x103),.w(w39_102),.acc(r39_102),.res(r39_103),.clk(clk),.wout(w39_103));
	PE pe39_104(.x(x104),.w(w39_103),.acc(r39_103),.res(r39_104),.clk(clk),.wout(w39_104));
	PE pe39_105(.x(x105),.w(w39_104),.acc(r39_104),.res(r39_105),.clk(clk),.wout(w39_105));
	PE pe39_106(.x(x106),.w(w39_105),.acc(r39_105),.res(r39_106),.clk(clk),.wout(w39_106));
	PE pe39_107(.x(x107),.w(w39_106),.acc(r39_106),.res(r39_107),.clk(clk),.wout(w39_107));
	PE pe39_108(.x(x108),.w(w39_107),.acc(r39_107),.res(r39_108),.clk(clk),.wout(w39_108));
	PE pe39_109(.x(x109),.w(w39_108),.acc(r39_108),.res(r39_109),.clk(clk),.wout(w39_109));
	PE pe39_110(.x(x110),.w(w39_109),.acc(r39_109),.res(r39_110),.clk(clk),.wout(w39_110));
	PE pe39_111(.x(x111),.w(w39_110),.acc(r39_110),.res(r39_111),.clk(clk),.wout(w39_111));
	PE pe39_112(.x(x112),.w(w39_111),.acc(r39_111),.res(r39_112),.clk(clk),.wout(w39_112));
	PE pe39_113(.x(x113),.w(w39_112),.acc(r39_112),.res(r39_113),.clk(clk),.wout(w39_113));
	PE pe39_114(.x(x114),.w(w39_113),.acc(r39_113),.res(r39_114),.clk(clk),.wout(w39_114));
	PE pe39_115(.x(x115),.w(w39_114),.acc(r39_114),.res(r39_115),.clk(clk),.wout(w39_115));
	PE pe39_116(.x(x116),.w(w39_115),.acc(r39_115),.res(r39_116),.clk(clk),.wout(w39_116));
	PE pe39_117(.x(x117),.w(w39_116),.acc(r39_116),.res(r39_117),.clk(clk),.wout(w39_117));
	PE pe39_118(.x(x118),.w(w39_117),.acc(r39_117),.res(r39_118),.clk(clk),.wout(w39_118));
	PE pe39_119(.x(x119),.w(w39_118),.acc(r39_118),.res(r39_119),.clk(clk),.wout(w39_119));
	PE pe39_120(.x(x120),.w(w39_119),.acc(r39_119),.res(r39_120),.clk(clk),.wout(w39_120));
	PE pe39_121(.x(x121),.w(w39_120),.acc(r39_120),.res(r39_121),.clk(clk),.wout(w39_121));
	PE pe39_122(.x(x122),.w(w39_121),.acc(r39_121),.res(r39_122),.clk(clk),.wout(w39_122));
	PE pe39_123(.x(x123),.w(w39_122),.acc(r39_122),.res(r39_123),.clk(clk),.wout(w39_123));
	PE pe39_124(.x(x124),.w(w39_123),.acc(r39_123),.res(r39_124),.clk(clk),.wout(w39_124));
	PE pe39_125(.x(x125),.w(w39_124),.acc(r39_124),.res(r39_125),.clk(clk),.wout(w39_125));
	PE pe39_126(.x(x126),.w(w39_125),.acc(r39_125),.res(r39_126),.clk(clk),.wout(w39_126));
	PE pe39_127(.x(x127),.w(w39_126),.acc(r39_126),.res(result39),.clk(clk),.wout(weight39));

	PE pe40_0(.x(x0),.w(w40),.acc(32'h0),.res(r40_0),.clk(clk),.wout(w40_0));
	PE pe40_1(.x(x1),.w(w40_0),.acc(r40_0),.res(r40_1),.clk(clk),.wout(w40_1));
	PE pe40_2(.x(x2),.w(w40_1),.acc(r40_1),.res(r40_2),.clk(clk),.wout(w40_2));
	PE pe40_3(.x(x3),.w(w40_2),.acc(r40_2),.res(r40_3),.clk(clk),.wout(w40_3));
	PE pe40_4(.x(x4),.w(w40_3),.acc(r40_3),.res(r40_4),.clk(clk),.wout(w40_4));
	PE pe40_5(.x(x5),.w(w40_4),.acc(r40_4),.res(r40_5),.clk(clk),.wout(w40_5));
	PE pe40_6(.x(x6),.w(w40_5),.acc(r40_5),.res(r40_6),.clk(clk),.wout(w40_6));
	PE pe40_7(.x(x7),.w(w40_6),.acc(r40_6),.res(r40_7),.clk(clk),.wout(w40_7));
	PE pe40_8(.x(x8),.w(w40_7),.acc(r40_7),.res(r40_8),.clk(clk),.wout(w40_8));
	PE pe40_9(.x(x9),.w(w40_8),.acc(r40_8),.res(r40_9),.clk(clk),.wout(w40_9));
	PE pe40_10(.x(x10),.w(w40_9),.acc(r40_9),.res(r40_10),.clk(clk),.wout(w40_10));
	PE pe40_11(.x(x11),.w(w40_10),.acc(r40_10),.res(r40_11),.clk(clk),.wout(w40_11));
	PE pe40_12(.x(x12),.w(w40_11),.acc(r40_11),.res(r40_12),.clk(clk),.wout(w40_12));
	PE pe40_13(.x(x13),.w(w40_12),.acc(r40_12),.res(r40_13),.clk(clk),.wout(w40_13));
	PE pe40_14(.x(x14),.w(w40_13),.acc(r40_13),.res(r40_14),.clk(clk),.wout(w40_14));
	PE pe40_15(.x(x15),.w(w40_14),.acc(r40_14),.res(r40_15),.clk(clk),.wout(w40_15));
	PE pe40_16(.x(x16),.w(w40_15),.acc(r40_15),.res(r40_16),.clk(clk),.wout(w40_16));
	PE pe40_17(.x(x17),.w(w40_16),.acc(r40_16),.res(r40_17),.clk(clk),.wout(w40_17));
	PE pe40_18(.x(x18),.w(w40_17),.acc(r40_17),.res(r40_18),.clk(clk),.wout(w40_18));
	PE pe40_19(.x(x19),.w(w40_18),.acc(r40_18),.res(r40_19),.clk(clk),.wout(w40_19));
	PE pe40_20(.x(x20),.w(w40_19),.acc(r40_19),.res(r40_20),.clk(clk),.wout(w40_20));
	PE pe40_21(.x(x21),.w(w40_20),.acc(r40_20),.res(r40_21),.clk(clk),.wout(w40_21));
	PE pe40_22(.x(x22),.w(w40_21),.acc(r40_21),.res(r40_22),.clk(clk),.wout(w40_22));
	PE pe40_23(.x(x23),.w(w40_22),.acc(r40_22),.res(r40_23),.clk(clk),.wout(w40_23));
	PE pe40_24(.x(x24),.w(w40_23),.acc(r40_23),.res(r40_24),.clk(clk),.wout(w40_24));
	PE pe40_25(.x(x25),.w(w40_24),.acc(r40_24),.res(r40_25),.clk(clk),.wout(w40_25));
	PE pe40_26(.x(x26),.w(w40_25),.acc(r40_25),.res(r40_26),.clk(clk),.wout(w40_26));
	PE pe40_27(.x(x27),.w(w40_26),.acc(r40_26),.res(r40_27),.clk(clk),.wout(w40_27));
	PE pe40_28(.x(x28),.w(w40_27),.acc(r40_27),.res(r40_28),.clk(clk),.wout(w40_28));
	PE pe40_29(.x(x29),.w(w40_28),.acc(r40_28),.res(r40_29),.clk(clk),.wout(w40_29));
	PE pe40_30(.x(x30),.w(w40_29),.acc(r40_29),.res(r40_30),.clk(clk),.wout(w40_30));
	PE pe40_31(.x(x31),.w(w40_30),.acc(r40_30),.res(r40_31),.clk(clk),.wout(w40_31));
	PE pe40_32(.x(x32),.w(w40_31),.acc(r40_31),.res(r40_32),.clk(clk),.wout(w40_32));
	PE pe40_33(.x(x33),.w(w40_32),.acc(r40_32),.res(r40_33),.clk(clk),.wout(w40_33));
	PE pe40_34(.x(x34),.w(w40_33),.acc(r40_33),.res(r40_34),.clk(clk),.wout(w40_34));
	PE pe40_35(.x(x35),.w(w40_34),.acc(r40_34),.res(r40_35),.clk(clk),.wout(w40_35));
	PE pe40_36(.x(x36),.w(w40_35),.acc(r40_35),.res(r40_36),.clk(clk),.wout(w40_36));
	PE pe40_37(.x(x37),.w(w40_36),.acc(r40_36),.res(r40_37),.clk(clk),.wout(w40_37));
	PE pe40_38(.x(x38),.w(w40_37),.acc(r40_37),.res(r40_38),.clk(clk),.wout(w40_38));
	PE pe40_39(.x(x39),.w(w40_38),.acc(r40_38),.res(r40_39),.clk(clk),.wout(w40_39));
	PE pe40_40(.x(x40),.w(w40_39),.acc(r40_39),.res(r40_40),.clk(clk),.wout(w40_40));
	PE pe40_41(.x(x41),.w(w40_40),.acc(r40_40),.res(r40_41),.clk(clk),.wout(w40_41));
	PE pe40_42(.x(x42),.w(w40_41),.acc(r40_41),.res(r40_42),.clk(clk),.wout(w40_42));
	PE pe40_43(.x(x43),.w(w40_42),.acc(r40_42),.res(r40_43),.clk(clk),.wout(w40_43));
	PE pe40_44(.x(x44),.w(w40_43),.acc(r40_43),.res(r40_44),.clk(clk),.wout(w40_44));
	PE pe40_45(.x(x45),.w(w40_44),.acc(r40_44),.res(r40_45),.clk(clk),.wout(w40_45));
	PE pe40_46(.x(x46),.w(w40_45),.acc(r40_45),.res(r40_46),.clk(clk),.wout(w40_46));
	PE pe40_47(.x(x47),.w(w40_46),.acc(r40_46),.res(r40_47),.clk(clk),.wout(w40_47));
	PE pe40_48(.x(x48),.w(w40_47),.acc(r40_47),.res(r40_48),.clk(clk),.wout(w40_48));
	PE pe40_49(.x(x49),.w(w40_48),.acc(r40_48),.res(r40_49),.clk(clk),.wout(w40_49));
	PE pe40_50(.x(x50),.w(w40_49),.acc(r40_49),.res(r40_50),.clk(clk),.wout(w40_50));
	PE pe40_51(.x(x51),.w(w40_50),.acc(r40_50),.res(r40_51),.clk(clk),.wout(w40_51));
	PE pe40_52(.x(x52),.w(w40_51),.acc(r40_51),.res(r40_52),.clk(clk),.wout(w40_52));
	PE pe40_53(.x(x53),.w(w40_52),.acc(r40_52),.res(r40_53),.clk(clk),.wout(w40_53));
	PE pe40_54(.x(x54),.w(w40_53),.acc(r40_53),.res(r40_54),.clk(clk),.wout(w40_54));
	PE pe40_55(.x(x55),.w(w40_54),.acc(r40_54),.res(r40_55),.clk(clk),.wout(w40_55));
	PE pe40_56(.x(x56),.w(w40_55),.acc(r40_55),.res(r40_56),.clk(clk),.wout(w40_56));
	PE pe40_57(.x(x57),.w(w40_56),.acc(r40_56),.res(r40_57),.clk(clk),.wout(w40_57));
	PE pe40_58(.x(x58),.w(w40_57),.acc(r40_57),.res(r40_58),.clk(clk),.wout(w40_58));
	PE pe40_59(.x(x59),.w(w40_58),.acc(r40_58),.res(r40_59),.clk(clk),.wout(w40_59));
	PE pe40_60(.x(x60),.w(w40_59),.acc(r40_59),.res(r40_60),.clk(clk),.wout(w40_60));
	PE pe40_61(.x(x61),.w(w40_60),.acc(r40_60),.res(r40_61),.clk(clk),.wout(w40_61));
	PE pe40_62(.x(x62),.w(w40_61),.acc(r40_61),.res(r40_62),.clk(clk),.wout(w40_62));
	PE pe40_63(.x(x63),.w(w40_62),.acc(r40_62),.res(r40_63),.clk(clk),.wout(w40_63));
	PE pe40_64(.x(x64),.w(w40_63),.acc(r40_63),.res(r40_64),.clk(clk),.wout(w40_64));
	PE pe40_65(.x(x65),.w(w40_64),.acc(r40_64),.res(r40_65),.clk(clk),.wout(w40_65));
	PE pe40_66(.x(x66),.w(w40_65),.acc(r40_65),.res(r40_66),.clk(clk),.wout(w40_66));
	PE pe40_67(.x(x67),.w(w40_66),.acc(r40_66),.res(r40_67),.clk(clk),.wout(w40_67));
	PE pe40_68(.x(x68),.w(w40_67),.acc(r40_67),.res(r40_68),.clk(clk),.wout(w40_68));
	PE pe40_69(.x(x69),.w(w40_68),.acc(r40_68),.res(r40_69),.clk(clk),.wout(w40_69));
	PE pe40_70(.x(x70),.w(w40_69),.acc(r40_69),.res(r40_70),.clk(clk),.wout(w40_70));
	PE pe40_71(.x(x71),.w(w40_70),.acc(r40_70),.res(r40_71),.clk(clk),.wout(w40_71));
	PE pe40_72(.x(x72),.w(w40_71),.acc(r40_71),.res(r40_72),.clk(clk),.wout(w40_72));
	PE pe40_73(.x(x73),.w(w40_72),.acc(r40_72),.res(r40_73),.clk(clk),.wout(w40_73));
	PE pe40_74(.x(x74),.w(w40_73),.acc(r40_73),.res(r40_74),.clk(clk),.wout(w40_74));
	PE pe40_75(.x(x75),.w(w40_74),.acc(r40_74),.res(r40_75),.clk(clk),.wout(w40_75));
	PE pe40_76(.x(x76),.w(w40_75),.acc(r40_75),.res(r40_76),.clk(clk),.wout(w40_76));
	PE pe40_77(.x(x77),.w(w40_76),.acc(r40_76),.res(r40_77),.clk(clk),.wout(w40_77));
	PE pe40_78(.x(x78),.w(w40_77),.acc(r40_77),.res(r40_78),.clk(clk),.wout(w40_78));
	PE pe40_79(.x(x79),.w(w40_78),.acc(r40_78),.res(r40_79),.clk(clk),.wout(w40_79));
	PE pe40_80(.x(x80),.w(w40_79),.acc(r40_79),.res(r40_80),.clk(clk),.wout(w40_80));
	PE pe40_81(.x(x81),.w(w40_80),.acc(r40_80),.res(r40_81),.clk(clk),.wout(w40_81));
	PE pe40_82(.x(x82),.w(w40_81),.acc(r40_81),.res(r40_82),.clk(clk),.wout(w40_82));
	PE pe40_83(.x(x83),.w(w40_82),.acc(r40_82),.res(r40_83),.clk(clk),.wout(w40_83));
	PE pe40_84(.x(x84),.w(w40_83),.acc(r40_83),.res(r40_84),.clk(clk),.wout(w40_84));
	PE pe40_85(.x(x85),.w(w40_84),.acc(r40_84),.res(r40_85),.clk(clk),.wout(w40_85));
	PE pe40_86(.x(x86),.w(w40_85),.acc(r40_85),.res(r40_86),.clk(clk),.wout(w40_86));
	PE pe40_87(.x(x87),.w(w40_86),.acc(r40_86),.res(r40_87),.clk(clk),.wout(w40_87));
	PE pe40_88(.x(x88),.w(w40_87),.acc(r40_87),.res(r40_88),.clk(clk),.wout(w40_88));
	PE pe40_89(.x(x89),.w(w40_88),.acc(r40_88),.res(r40_89),.clk(clk),.wout(w40_89));
	PE pe40_90(.x(x90),.w(w40_89),.acc(r40_89),.res(r40_90),.clk(clk),.wout(w40_90));
	PE pe40_91(.x(x91),.w(w40_90),.acc(r40_90),.res(r40_91),.clk(clk),.wout(w40_91));
	PE pe40_92(.x(x92),.w(w40_91),.acc(r40_91),.res(r40_92),.clk(clk),.wout(w40_92));
	PE pe40_93(.x(x93),.w(w40_92),.acc(r40_92),.res(r40_93),.clk(clk),.wout(w40_93));
	PE pe40_94(.x(x94),.w(w40_93),.acc(r40_93),.res(r40_94),.clk(clk),.wout(w40_94));
	PE pe40_95(.x(x95),.w(w40_94),.acc(r40_94),.res(r40_95),.clk(clk),.wout(w40_95));
	PE pe40_96(.x(x96),.w(w40_95),.acc(r40_95),.res(r40_96),.clk(clk),.wout(w40_96));
	PE pe40_97(.x(x97),.w(w40_96),.acc(r40_96),.res(r40_97),.clk(clk),.wout(w40_97));
	PE pe40_98(.x(x98),.w(w40_97),.acc(r40_97),.res(r40_98),.clk(clk),.wout(w40_98));
	PE pe40_99(.x(x99),.w(w40_98),.acc(r40_98),.res(r40_99),.clk(clk),.wout(w40_99));
	PE pe40_100(.x(x100),.w(w40_99),.acc(r40_99),.res(r40_100),.clk(clk),.wout(w40_100));
	PE pe40_101(.x(x101),.w(w40_100),.acc(r40_100),.res(r40_101),.clk(clk),.wout(w40_101));
	PE pe40_102(.x(x102),.w(w40_101),.acc(r40_101),.res(r40_102),.clk(clk),.wout(w40_102));
	PE pe40_103(.x(x103),.w(w40_102),.acc(r40_102),.res(r40_103),.clk(clk),.wout(w40_103));
	PE pe40_104(.x(x104),.w(w40_103),.acc(r40_103),.res(r40_104),.clk(clk),.wout(w40_104));
	PE pe40_105(.x(x105),.w(w40_104),.acc(r40_104),.res(r40_105),.clk(clk),.wout(w40_105));
	PE pe40_106(.x(x106),.w(w40_105),.acc(r40_105),.res(r40_106),.clk(clk),.wout(w40_106));
	PE pe40_107(.x(x107),.w(w40_106),.acc(r40_106),.res(r40_107),.clk(clk),.wout(w40_107));
	PE pe40_108(.x(x108),.w(w40_107),.acc(r40_107),.res(r40_108),.clk(clk),.wout(w40_108));
	PE pe40_109(.x(x109),.w(w40_108),.acc(r40_108),.res(r40_109),.clk(clk),.wout(w40_109));
	PE pe40_110(.x(x110),.w(w40_109),.acc(r40_109),.res(r40_110),.clk(clk),.wout(w40_110));
	PE pe40_111(.x(x111),.w(w40_110),.acc(r40_110),.res(r40_111),.clk(clk),.wout(w40_111));
	PE pe40_112(.x(x112),.w(w40_111),.acc(r40_111),.res(r40_112),.clk(clk),.wout(w40_112));
	PE pe40_113(.x(x113),.w(w40_112),.acc(r40_112),.res(r40_113),.clk(clk),.wout(w40_113));
	PE pe40_114(.x(x114),.w(w40_113),.acc(r40_113),.res(r40_114),.clk(clk),.wout(w40_114));
	PE pe40_115(.x(x115),.w(w40_114),.acc(r40_114),.res(r40_115),.clk(clk),.wout(w40_115));
	PE pe40_116(.x(x116),.w(w40_115),.acc(r40_115),.res(r40_116),.clk(clk),.wout(w40_116));
	PE pe40_117(.x(x117),.w(w40_116),.acc(r40_116),.res(r40_117),.clk(clk),.wout(w40_117));
	PE pe40_118(.x(x118),.w(w40_117),.acc(r40_117),.res(r40_118),.clk(clk),.wout(w40_118));
	PE pe40_119(.x(x119),.w(w40_118),.acc(r40_118),.res(r40_119),.clk(clk),.wout(w40_119));
	PE pe40_120(.x(x120),.w(w40_119),.acc(r40_119),.res(r40_120),.clk(clk),.wout(w40_120));
	PE pe40_121(.x(x121),.w(w40_120),.acc(r40_120),.res(r40_121),.clk(clk),.wout(w40_121));
	PE pe40_122(.x(x122),.w(w40_121),.acc(r40_121),.res(r40_122),.clk(clk),.wout(w40_122));
	PE pe40_123(.x(x123),.w(w40_122),.acc(r40_122),.res(r40_123),.clk(clk),.wout(w40_123));
	PE pe40_124(.x(x124),.w(w40_123),.acc(r40_123),.res(r40_124),.clk(clk),.wout(w40_124));
	PE pe40_125(.x(x125),.w(w40_124),.acc(r40_124),.res(r40_125),.clk(clk),.wout(w40_125));
	PE pe40_126(.x(x126),.w(w40_125),.acc(r40_125),.res(r40_126),.clk(clk),.wout(w40_126));
	PE pe40_127(.x(x127),.w(w40_126),.acc(r40_126),.res(result40),.clk(clk),.wout(weight40));

	PE pe41_0(.x(x0),.w(w41),.acc(32'h0),.res(r41_0),.clk(clk),.wout(w41_0));
	PE pe41_1(.x(x1),.w(w41_0),.acc(r41_0),.res(r41_1),.clk(clk),.wout(w41_1));
	PE pe41_2(.x(x2),.w(w41_1),.acc(r41_1),.res(r41_2),.clk(clk),.wout(w41_2));
	PE pe41_3(.x(x3),.w(w41_2),.acc(r41_2),.res(r41_3),.clk(clk),.wout(w41_3));
	PE pe41_4(.x(x4),.w(w41_3),.acc(r41_3),.res(r41_4),.clk(clk),.wout(w41_4));
	PE pe41_5(.x(x5),.w(w41_4),.acc(r41_4),.res(r41_5),.clk(clk),.wout(w41_5));
	PE pe41_6(.x(x6),.w(w41_5),.acc(r41_5),.res(r41_6),.clk(clk),.wout(w41_6));
	PE pe41_7(.x(x7),.w(w41_6),.acc(r41_6),.res(r41_7),.clk(clk),.wout(w41_7));
	PE pe41_8(.x(x8),.w(w41_7),.acc(r41_7),.res(r41_8),.clk(clk),.wout(w41_8));
	PE pe41_9(.x(x9),.w(w41_8),.acc(r41_8),.res(r41_9),.clk(clk),.wout(w41_9));
	PE pe41_10(.x(x10),.w(w41_9),.acc(r41_9),.res(r41_10),.clk(clk),.wout(w41_10));
	PE pe41_11(.x(x11),.w(w41_10),.acc(r41_10),.res(r41_11),.clk(clk),.wout(w41_11));
	PE pe41_12(.x(x12),.w(w41_11),.acc(r41_11),.res(r41_12),.clk(clk),.wout(w41_12));
	PE pe41_13(.x(x13),.w(w41_12),.acc(r41_12),.res(r41_13),.clk(clk),.wout(w41_13));
	PE pe41_14(.x(x14),.w(w41_13),.acc(r41_13),.res(r41_14),.clk(clk),.wout(w41_14));
	PE pe41_15(.x(x15),.w(w41_14),.acc(r41_14),.res(r41_15),.clk(clk),.wout(w41_15));
	PE pe41_16(.x(x16),.w(w41_15),.acc(r41_15),.res(r41_16),.clk(clk),.wout(w41_16));
	PE pe41_17(.x(x17),.w(w41_16),.acc(r41_16),.res(r41_17),.clk(clk),.wout(w41_17));
	PE pe41_18(.x(x18),.w(w41_17),.acc(r41_17),.res(r41_18),.clk(clk),.wout(w41_18));
	PE pe41_19(.x(x19),.w(w41_18),.acc(r41_18),.res(r41_19),.clk(clk),.wout(w41_19));
	PE pe41_20(.x(x20),.w(w41_19),.acc(r41_19),.res(r41_20),.clk(clk),.wout(w41_20));
	PE pe41_21(.x(x21),.w(w41_20),.acc(r41_20),.res(r41_21),.clk(clk),.wout(w41_21));
	PE pe41_22(.x(x22),.w(w41_21),.acc(r41_21),.res(r41_22),.clk(clk),.wout(w41_22));
	PE pe41_23(.x(x23),.w(w41_22),.acc(r41_22),.res(r41_23),.clk(clk),.wout(w41_23));
	PE pe41_24(.x(x24),.w(w41_23),.acc(r41_23),.res(r41_24),.clk(clk),.wout(w41_24));
	PE pe41_25(.x(x25),.w(w41_24),.acc(r41_24),.res(r41_25),.clk(clk),.wout(w41_25));
	PE pe41_26(.x(x26),.w(w41_25),.acc(r41_25),.res(r41_26),.clk(clk),.wout(w41_26));
	PE pe41_27(.x(x27),.w(w41_26),.acc(r41_26),.res(r41_27),.clk(clk),.wout(w41_27));
	PE pe41_28(.x(x28),.w(w41_27),.acc(r41_27),.res(r41_28),.clk(clk),.wout(w41_28));
	PE pe41_29(.x(x29),.w(w41_28),.acc(r41_28),.res(r41_29),.clk(clk),.wout(w41_29));
	PE pe41_30(.x(x30),.w(w41_29),.acc(r41_29),.res(r41_30),.clk(clk),.wout(w41_30));
	PE pe41_31(.x(x31),.w(w41_30),.acc(r41_30),.res(r41_31),.clk(clk),.wout(w41_31));
	PE pe41_32(.x(x32),.w(w41_31),.acc(r41_31),.res(r41_32),.clk(clk),.wout(w41_32));
	PE pe41_33(.x(x33),.w(w41_32),.acc(r41_32),.res(r41_33),.clk(clk),.wout(w41_33));
	PE pe41_34(.x(x34),.w(w41_33),.acc(r41_33),.res(r41_34),.clk(clk),.wout(w41_34));
	PE pe41_35(.x(x35),.w(w41_34),.acc(r41_34),.res(r41_35),.clk(clk),.wout(w41_35));
	PE pe41_36(.x(x36),.w(w41_35),.acc(r41_35),.res(r41_36),.clk(clk),.wout(w41_36));
	PE pe41_37(.x(x37),.w(w41_36),.acc(r41_36),.res(r41_37),.clk(clk),.wout(w41_37));
	PE pe41_38(.x(x38),.w(w41_37),.acc(r41_37),.res(r41_38),.clk(clk),.wout(w41_38));
	PE pe41_39(.x(x39),.w(w41_38),.acc(r41_38),.res(r41_39),.clk(clk),.wout(w41_39));
	PE pe41_40(.x(x40),.w(w41_39),.acc(r41_39),.res(r41_40),.clk(clk),.wout(w41_40));
	PE pe41_41(.x(x41),.w(w41_40),.acc(r41_40),.res(r41_41),.clk(clk),.wout(w41_41));
	PE pe41_42(.x(x42),.w(w41_41),.acc(r41_41),.res(r41_42),.clk(clk),.wout(w41_42));
	PE pe41_43(.x(x43),.w(w41_42),.acc(r41_42),.res(r41_43),.clk(clk),.wout(w41_43));
	PE pe41_44(.x(x44),.w(w41_43),.acc(r41_43),.res(r41_44),.clk(clk),.wout(w41_44));
	PE pe41_45(.x(x45),.w(w41_44),.acc(r41_44),.res(r41_45),.clk(clk),.wout(w41_45));
	PE pe41_46(.x(x46),.w(w41_45),.acc(r41_45),.res(r41_46),.clk(clk),.wout(w41_46));
	PE pe41_47(.x(x47),.w(w41_46),.acc(r41_46),.res(r41_47),.clk(clk),.wout(w41_47));
	PE pe41_48(.x(x48),.w(w41_47),.acc(r41_47),.res(r41_48),.clk(clk),.wout(w41_48));
	PE pe41_49(.x(x49),.w(w41_48),.acc(r41_48),.res(r41_49),.clk(clk),.wout(w41_49));
	PE pe41_50(.x(x50),.w(w41_49),.acc(r41_49),.res(r41_50),.clk(clk),.wout(w41_50));
	PE pe41_51(.x(x51),.w(w41_50),.acc(r41_50),.res(r41_51),.clk(clk),.wout(w41_51));
	PE pe41_52(.x(x52),.w(w41_51),.acc(r41_51),.res(r41_52),.clk(clk),.wout(w41_52));
	PE pe41_53(.x(x53),.w(w41_52),.acc(r41_52),.res(r41_53),.clk(clk),.wout(w41_53));
	PE pe41_54(.x(x54),.w(w41_53),.acc(r41_53),.res(r41_54),.clk(clk),.wout(w41_54));
	PE pe41_55(.x(x55),.w(w41_54),.acc(r41_54),.res(r41_55),.clk(clk),.wout(w41_55));
	PE pe41_56(.x(x56),.w(w41_55),.acc(r41_55),.res(r41_56),.clk(clk),.wout(w41_56));
	PE pe41_57(.x(x57),.w(w41_56),.acc(r41_56),.res(r41_57),.clk(clk),.wout(w41_57));
	PE pe41_58(.x(x58),.w(w41_57),.acc(r41_57),.res(r41_58),.clk(clk),.wout(w41_58));
	PE pe41_59(.x(x59),.w(w41_58),.acc(r41_58),.res(r41_59),.clk(clk),.wout(w41_59));
	PE pe41_60(.x(x60),.w(w41_59),.acc(r41_59),.res(r41_60),.clk(clk),.wout(w41_60));
	PE pe41_61(.x(x61),.w(w41_60),.acc(r41_60),.res(r41_61),.clk(clk),.wout(w41_61));
	PE pe41_62(.x(x62),.w(w41_61),.acc(r41_61),.res(r41_62),.clk(clk),.wout(w41_62));
	PE pe41_63(.x(x63),.w(w41_62),.acc(r41_62),.res(r41_63),.clk(clk),.wout(w41_63));
	PE pe41_64(.x(x64),.w(w41_63),.acc(r41_63),.res(r41_64),.clk(clk),.wout(w41_64));
	PE pe41_65(.x(x65),.w(w41_64),.acc(r41_64),.res(r41_65),.clk(clk),.wout(w41_65));
	PE pe41_66(.x(x66),.w(w41_65),.acc(r41_65),.res(r41_66),.clk(clk),.wout(w41_66));
	PE pe41_67(.x(x67),.w(w41_66),.acc(r41_66),.res(r41_67),.clk(clk),.wout(w41_67));
	PE pe41_68(.x(x68),.w(w41_67),.acc(r41_67),.res(r41_68),.clk(clk),.wout(w41_68));
	PE pe41_69(.x(x69),.w(w41_68),.acc(r41_68),.res(r41_69),.clk(clk),.wout(w41_69));
	PE pe41_70(.x(x70),.w(w41_69),.acc(r41_69),.res(r41_70),.clk(clk),.wout(w41_70));
	PE pe41_71(.x(x71),.w(w41_70),.acc(r41_70),.res(r41_71),.clk(clk),.wout(w41_71));
	PE pe41_72(.x(x72),.w(w41_71),.acc(r41_71),.res(r41_72),.clk(clk),.wout(w41_72));
	PE pe41_73(.x(x73),.w(w41_72),.acc(r41_72),.res(r41_73),.clk(clk),.wout(w41_73));
	PE pe41_74(.x(x74),.w(w41_73),.acc(r41_73),.res(r41_74),.clk(clk),.wout(w41_74));
	PE pe41_75(.x(x75),.w(w41_74),.acc(r41_74),.res(r41_75),.clk(clk),.wout(w41_75));
	PE pe41_76(.x(x76),.w(w41_75),.acc(r41_75),.res(r41_76),.clk(clk),.wout(w41_76));
	PE pe41_77(.x(x77),.w(w41_76),.acc(r41_76),.res(r41_77),.clk(clk),.wout(w41_77));
	PE pe41_78(.x(x78),.w(w41_77),.acc(r41_77),.res(r41_78),.clk(clk),.wout(w41_78));
	PE pe41_79(.x(x79),.w(w41_78),.acc(r41_78),.res(r41_79),.clk(clk),.wout(w41_79));
	PE pe41_80(.x(x80),.w(w41_79),.acc(r41_79),.res(r41_80),.clk(clk),.wout(w41_80));
	PE pe41_81(.x(x81),.w(w41_80),.acc(r41_80),.res(r41_81),.clk(clk),.wout(w41_81));
	PE pe41_82(.x(x82),.w(w41_81),.acc(r41_81),.res(r41_82),.clk(clk),.wout(w41_82));
	PE pe41_83(.x(x83),.w(w41_82),.acc(r41_82),.res(r41_83),.clk(clk),.wout(w41_83));
	PE pe41_84(.x(x84),.w(w41_83),.acc(r41_83),.res(r41_84),.clk(clk),.wout(w41_84));
	PE pe41_85(.x(x85),.w(w41_84),.acc(r41_84),.res(r41_85),.clk(clk),.wout(w41_85));
	PE pe41_86(.x(x86),.w(w41_85),.acc(r41_85),.res(r41_86),.clk(clk),.wout(w41_86));
	PE pe41_87(.x(x87),.w(w41_86),.acc(r41_86),.res(r41_87),.clk(clk),.wout(w41_87));
	PE pe41_88(.x(x88),.w(w41_87),.acc(r41_87),.res(r41_88),.clk(clk),.wout(w41_88));
	PE pe41_89(.x(x89),.w(w41_88),.acc(r41_88),.res(r41_89),.clk(clk),.wout(w41_89));
	PE pe41_90(.x(x90),.w(w41_89),.acc(r41_89),.res(r41_90),.clk(clk),.wout(w41_90));
	PE pe41_91(.x(x91),.w(w41_90),.acc(r41_90),.res(r41_91),.clk(clk),.wout(w41_91));
	PE pe41_92(.x(x92),.w(w41_91),.acc(r41_91),.res(r41_92),.clk(clk),.wout(w41_92));
	PE pe41_93(.x(x93),.w(w41_92),.acc(r41_92),.res(r41_93),.clk(clk),.wout(w41_93));
	PE pe41_94(.x(x94),.w(w41_93),.acc(r41_93),.res(r41_94),.clk(clk),.wout(w41_94));
	PE pe41_95(.x(x95),.w(w41_94),.acc(r41_94),.res(r41_95),.clk(clk),.wout(w41_95));
	PE pe41_96(.x(x96),.w(w41_95),.acc(r41_95),.res(r41_96),.clk(clk),.wout(w41_96));
	PE pe41_97(.x(x97),.w(w41_96),.acc(r41_96),.res(r41_97),.clk(clk),.wout(w41_97));
	PE pe41_98(.x(x98),.w(w41_97),.acc(r41_97),.res(r41_98),.clk(clk),.wout(w41_98));
	PE pe41_99(.x(x99),.w(w41_98),.acc(r41_98),.res(r41_99),.clk(clk),.wout(w41_99));
	PE pe41_100(.x(x100),.w(w41_99),.acc(r41_99),.res(r41_100),.clk(clk),.wout(w41_100));
	PE pe41_101(.x(x101),.w(w41_100),.acc(r41_100),.res(r41_101),.clk(clk),.wout(w41_101));
	PE pe41_102(.x(x102),.w(w41_101),.acc(r41_101),.res(r41_102),.clk(clk),.wout(w41_102));
	PE pe41_103(.x(x103),.w(w41_102),.acc(r41_102),.res(r41_103),.clk(clk),.wout(w41_103));
	PE pe41_104(.x(x104),.w(w41_103),.acc(r41_103),.res(r41_104),.clk(clk),.wout(w41_104));
	PE pe41_105(.x(x105),.w(w41_104),.acc(r41_104),.res(r41_105),.clk(clk),.wout(w41_105));
	PE pe41_106(.x(x106),.w(w41_105),.acc(r41_105),.res(r41_106),.clk(clk),.wout(w41_106));
	PE pe41_107(.x(x107),.w(w41_106),.acc(r41_106),.res(r41_107),.clk(clk),.wout(w41_107));
	PE pe41_108(.x(x108),.w(w41_107),.acc(r41_107),.res(r41_108),.clk(clk),.wout(w41_108));
	PE pe41_109(.x(x109),.w(w41_108),.acc(r41_108),.res(r41_109),.clk(clk),.wout(w41_109));
	PE pe41_110(.x(x110),.w(w41_109),.acc(r41_109),.res(r41_110),.clk(clk),.wout(w41_110));
	PE pe41_111(.x(x111),.w(w41_110),.acc(r41_110),.res(r41_111),.clk(clk),.wout(w41_111));
	PE pe41_112(.x(x112),.w(w41_111),.acc(r41_111),.res(r41_112),.clk(clk),.wout(w41_112));
	PE pe41_113(.x(x113),.w(w41_112),.acc(r41_112),.res(r41_113),.clk(clk),.wout(w41_113));
	PE pe41_114(.x(x114),.w(w41_113),.acc(r41_113),.res(r41_114),.clk(clk),.wout(w41_114));
	PE pe41_115(.x(x115),.w(w41_114),.acc(r41_114),.res(r41_115),.clk(clk),.wout(w41_115));
	PE pe41_116(.x(x116),.w(w41_115),.acc(r41_115),.res(r41_116),.clk(clk),.wout(w41_116));
	PE pe41_117(.x(x117),.w(w41_116),.acc(r41_116),.res(r41_117),.clk(clk),.wout(w41_117));
	PE pe41_118(.x(x118),.w(w41_117),.acc(r41_117),.res(r41_118),.clk(clk),.wout(w41_118));
	PE pe41_119(.x(x119),.w(w41_118),.acc(r41_118),.res(r41_119),.clk(clk),.wout(w41_119));
	PE pe41_120(.x(x120),.w(w41_119),.acc(r41_119),.res(r41_120),.clk(clk),.wout(w41_120));
	PE pe41_121(.x(x121),.w(w41_120),.acc(r41_120),.res(r41_121),.clk(clk),.wout(w41_121));
	PE pe41_122(.x(x122),.w(w41_121),.acc(r41_121),.res(r41_122),.clk(clk),.wout(w41_122));
	PE pe41_123(.x(x123),.w(w41_122),.acc(r41_122),.res(r41_123),.clk(clk),.wout(w41_123));
	PE pe41_124(.x(x124),.w(w41_123),.acc(r41_123),.res(r41_124),.clk(clk),.wout(w41_124));
	PE pe41_125(.x(x125),.w(w41_124),.acc(r41_124),.res(r41_125),.clk(clk),.wout(w41_125));
	PE pe41_126(.x(x126),.w(w41_125),.acc(r41_125),.res(r41_126),.clk(clk),.wout(w41_126));
	PE pe41_127(.x(x127),.w(w41_126),.acc(r41_126),.res(result41),.clk(clk),.wout(weight41));

	PE pe42_0(.x(x0),.w(w42),.acc(32'h0),.res(r42_0),.clk(clk),.wout(w42_0));
	PE pe42_1(.x(x1),.w(w42_0),.acc(r42_0),.res(r42_1),.clk(clk),.wout(w42_1));
	PE pe42_2(.x(x2),.w(w42_1),.acc(r42_1),.res(r42_2),.clk(clk),.wout(w42_2));
	PE pe42_3(.x(x3),.w(w42_2),.acc(r42_2),.res(r42_3),.clk(clk),.wout(w42_3));
	PE pe42_4(.x(x4),.w(w42_3),.acc(r42_3),.res(r42_4),.clk(clk),.wout(w42_4));
	PE pe42_5(.x(x5),.w(w42_4),.acc(r42_4),.res(r42_5),.clk(clk),.wout(w42_5));
	PE pe42_6(.x(x6),.w(w42_5),.acc(r42_5),.res(r42_6),.clk(clk),.wout(w42_6));
	PE pe42_7(.x(x7),.w(w42_6),.acc(r42_6),.res(r42_7),.clk(clk),.wout(w42_7));
	PE pe42_8(.x(x8),.w(w42_7),.acc(r42_7),.res(r42_8),.clk(clk),.wout(w42_8));
	PE pe42_9(.x(x9),.w(w42_8),.acc(r42_8),.res(r42_9),.clk(clk),.wout(w42_9));
	PE pe42_10(.x(x10),.w(w42_9),.acc(r42_9),.res(r42_10),.clk(clk),.wout(w42_10));
	PE pe42_11(.x(x11),.w(w42_10),.acc(r42_10),.res(r42_11),.clk(clk),.wout(w42_11));
	PE pe42_12(.x(x12),.w(w42_11),.acc(r42_11),.res(r42_12),.clk(clk),.wout(w42_12));
	PE pe42_13(.x(x13),.w(w42_12),.acc(r42_12),.res(r42_13),.clk(clk),.wout(w42_13));
	PE pe42_14(.x(x14),.w(w42_13),.acc(r42_13),.res(r42_14),.clk(clk),.wout(w42_14));
	PE pe42_15(.x(x15),.w(w42_14),.acc(r42_14),.res(r42_15),.clk(clk),.wout(w42_15));
	PE pe42_16(.x(x16),.w(w42_15),.acc(r42_15),.res(r42_16),.clk(clk),.wout(w42_16));
	PE pe42_17(.x(x17),.w(w42_16),.acc(r42_16),.res(r42_17),.clk(clk),.wout(w42_17));
	PE pe42_18(.x(x18),.w(w42_17),.acc(r42_17),.res(r42_18),.clk(clk),.wout(w42_18));
	PE pe42_19(.x(x19),.w(w42_18),.acc(r42_18),.res(r42_19),.clk(clk),.wout(w42_19));
	PE pe42_20(.x(x20),.w(w42_19),.acc(r42_19),.res(r42_20),.clk(clk),.wout(w42_20));
	PE pe42_21(.x(x21),.w(w42_20),.acc(r42_20),.res(r42_21),.clk(clk),.wout(w42_21));
	PE pe42_22(.x(x22),.w(w42_21),.acc(r42_21),.res(r42_22),.clk(clk),.wout(w42_22));
	PE pe42_23(.x(x23),.w(w42_22),.acc(r42_22),.res(r42_23),.clk(clk),.wout(w42_23));
	PE pe42_24(.x(x24),.w(w42_23),.acc(r42_23),.res(r42_24),.clk(clk),.wout(w42_24));
	PE pe42_25(.x(x25),.w(w42_24),.acc(r42_24),.res(r42_25),.clk(clk),.wout(w42_25));
	PE pe42_26(.x(x26),.w(w42_25),.acc(r42_25),.res(r42_26),.clk(clk),.wout(w42_26));
	PE pe42_27(.x(x27),.w(w42_26),.acc(r42_26),.res(r42_27),.clk(clk),.wout(w42_27));
	PE pe42_28(.x(x28),.w(w42_27),.acc(r42_27),.res(r42_28),.clk(clk),.wout(w42_28));
	PE pe42_29(.x(x29),.w(w42_28),.acc(r42_28),.res(r42_29),.clk(clk),.wout(w42_29));
	PE pe42_30(.x(x30),.w(w42_29),.acc(r42_29),.res(r42_30),.clk(clk),.wout(w42_30));
	PE pe42_31(.x(x31),.w(w42_30),.acc(r42_30),.res(r42_31),.clk(clk),.wout(w42_31));
	PE pe42_32(.x(x32),.w(w42_31),.acc(r42_31),.res(r42_32),.clk(clk),.wout(w42_32));
	PE pe42_33(.x(x33),.w(w42_32),.acc(r42_32),.res(r42_33),.clk(clk),.wout(w42_33));
	PE pe42_34(.x(x34),.w(w42_33),.acc(r42_33),.res(r42_34),.clk(clk),.wout(w42_34));
	PE pe42_35(.x(x35),.w(w42_34),.acc(r42_34),.res(r42_35),.clk(clk),.wout(w42_35));
	PE pe42_36(.x(x36),.w(w42_35),.acc(r42_35),.res(r42_36),.clk(clk),.wout(w42_36));
	PE pe42_37(.x(x37),.w(w42_36),.acc(r42_36),.res(r42_37),.clk(clk),.wout(w42_37));
	PE pe42_38(.x(x38),.w(w42_37),.acc(r42_37),.res(r42_38),.clk(clk),.wout(w42_38));
	PE pe42_39(.x(x39),.w(w42_38),.acc(r42_38),.res(r42_39),.clk(clk),.wout(w42_39));
	PE pe42_40(.x(x40),.w(w42_39),.acc(r42_39),.res(r42_40),.clk(clk),.wout(w42_40));
	PE pe42_41(.x(x41),.w(w42_40),.acc(r42_40),.res(r42_41),.clk(clk),.wout(w42_41));
	PE pe42_42(.x(x42),.w(w42_41),.acc(r42_41),.res(r42_42),.clk(clk),.wout(w42_42));
	PE pe42_43(.x(x43),.w(w42_42),.acc(r42_42),.res(r42_43),.clk(clk),.wout(w42_43));
	PE pe42_44(.x(x44),.w(w42_43),.acc(r42_43),.res(r42_44),.clk(clk),.wout(w42_44));
	PE pe42_45(.x(x45),.w(w42_44),.acc(r42_44),.res(r42_45),.clk(clk),.wout(w42_45));
	PE pe42_46(.x(x46),.w(w42_45),.acc(r42_45),.res(r42_46),.clk(clk),.wout(w42_46));
	PE pe42_47(.x(x47),.w(w42_46),.acc(r42_46),.res(r42_47),.clk(clk),.wout(w42_47));
	PE pe42_48(.x(x48),.w(w42_47),.acc(r42_47),.res(r42_48),.clk(clk),.wout(w42_48));
	PE pe42_49(.x(x49),.w(w42_48),.acc(r42_48),.res(r42_49),.clk(clk),.wout(w42_49));
	PE pe42_50(.x(x50),.w(w42_49),.acc(r42_49),.res(r42_50),.clk(clk),.wout(w42_50));
	PE pe42_51(.x(x51),.w(w42_50),.acc(r42_50),.res(r42_51),.clk(clk),.wout(w42_51));
	PE pe42_52(.x(x52),.w(w42_51),.acc(r42_51),.res(r42_52),.clk(clk),.wout(w42_52));
	PE pe42_53(.x(x53),.w(w42_52),.acc(r42_52),.res(r42_53),.clk(clk),.wout(w42_53));
	PE pe42_54(.x(x54),.w(w42_53),.acc(r42_53),.res(r42_54),.clk(clk),.wout(w42_54));
	PE pe42_55(.x(x55),.w(w42_54),.acc(r42_54),.res(r42_55),.clk(clk),.wout(w42_55));
	PE pe42_56(.x(x56),.w(w42_55),.acc(r42_55),.res(r42_56),.clk(clk),.wout(w42_56));
	PE pe42_57(.x(x57),.w(w42_56),.acc(r42_56),.res(r42_57),.clk(clk),.wout(w42_57));
	PE pe42_58(.x(x58),.w(w42_57),.acc(r42_57),.res(r42_58),.clk(clk),.wout(w42_58));
	PE pe42_59(.x(x59),.w(w42_58),.acc(r42_58),.res(r42_59),.clk(clk),.wout(w42_59));
	PE pe42_60(.x(x60),.w(w42_59),.acc(r42_59),.res(r42_60),.clk(clk),.wout(w42_60));
	PE pe42_61(.x(x61),.w(w42_60),.acc(r42_60),.res(r42_61),.clk(clk),.wout(w42_61));
	PE pe42_62(.x(x62),.w(w42_61),.acc(r42_61),.res(r42_62),.clk(clk),.wout(w42_62));
	PE pe42_63(.x(x63),.w(w42_62),.acc(r42_62),.res(r42_63),.clk(clk),.wout(w42_63));
	PE pe42_64(.x(x64),.w(w42_63),.acc(r42_63),.res(r42_64),.clk(clk),.wout(w42_64));
	PE pe42_65(.x(x65),.w(w42_64),.acc(r42_64),.res(r42_65),.clk(clk),.wout(w42_65));
	PE pe42_66(.x(x66),.w(w42_65),.acc(r42_65),.res(r42_66),.clk(clk),.wout(w42_66));
	PE pe42_67(.x(x67),.w(w42_66),.acc(r42_66),.res(r42_67),.clk(clk),.wout(w42_67));
	PE pe42_68(.x(x68),.w(w42_67),.acc(r42_67),.res(r42_68),.clk(clk),.wout(w42_68));
	PE pe42_69(.x(x69),.w(w42_68),.acc(r42_68),.res(r42_69),.clk(clk),.wout(w42_69));
	PE pe42_70(.x(x70),.w(w42_69),.acc(r42_69),.res(r42_70),.clk(clk),.wout(w42_70));
	PE pe42_71(.x(x71),.w(w42_70),.acc(r42_70),.res(r42_71),.clk(clk),.wout(w42_71));
	PE pe42_72(.x(x72),.w(w42_71),.acc(r42_71),.res(r42_72),.clk(clk),.wout(w42_72));
	PE pe42_73(.x(x73),.w(w42_72),.acc(r42_72),.res(r42_73),.clk(clk),.wout(w42_73));
	PE pe42_74(.x(x74),.w(w42_73),.acc(r42_73),.res(r42_74),.clk(clk),.wout(w42_74));
	PE pe42_75(.x(x75),.w(w42_74),.acc(r42_74),.res(r42_75),.clk(clk),.wout(w42_75));
	PE pe42_76(.x(x76),.w(w42_75),.acc(r42_75),.res(r42_76),.clk(clk),.wout(w42_76));
	PE pe42_77(.x(x77),.w(w42_76),.acc(r42_76),.res(r42_77),.clk(clk),.wout(w42_77));
	PE pe42_78(.x(x78),.w(w42_77),.acc(r42_77),.res(r42_78),.clk(clk),.wout(w42_78));
	PE pe42_79(.x(x79),.w(w42_78),.acc(r42_78),.res(r42_79),.clk(clk),.wout(w42_79));
	PE pe42_80(.x(x80),.w(w42_79),.acc(r42_79),.res(r42_80),.clk(clk),.wout(w42_80));
	PE pe42_81(.x(x81),.w(w42_80),.acc(r42_80),.res(r42_81),.clk(clk),.wout(w42_81));
	PE pe42_82(.x(x82),.w(w42_81),.acc(r42_81),.res(r42_82),.clk(clk),.wout(w42_82));
	PE pe42_83(.x(x83),.w(w42_82),.acc(r42_82),.res(r42_83),.clk(clk),.wout(w42_83));
	PE pe42_84(.x(x84),.w(w42_83),.acc(r42_83),.res(r42_84),.clk(clk),.wout(w42_84));
	PE pe42_85(.x(x85),.w(w42_84),.acc(r42_84),.res(r42_85),.clk(clk),.wout(w42_85));
	PE pe42_86(.x(x86),.w(w42_85),.acc(r42_85),.res(r42_86),.clk(clk),.wout(w42_86));
	PE pe42_87(.x(x87),.w(w42_86),.acc(r42_86),.res(r42_87),.clk(clk),.wout(w42_87));
	PE pe42_88(.x(x88),.w(w42_87),.acc(r42_87),.res(r42_88),.clk(clk),.wout(w42_88));
	PE pe42_89(.x(x89),.w(w42_88),.acc(r42_88),.res(r42_89),.clk(clk),.wout(w42_89));
	PE pe42_90(.x(x90),.w(w42_89),.acc(r42_89),.res(r42_90),.clk(clk),.wout(w42_90));
	PE pe42_91(.x(x91),.w(w42_90),.acc(r42_90),.res(r42_91),.clk(clk),.wout(w42_91));
	PE pe42_92(.x(x92),.w(w42_91),.acc(r42_91),.res(r42_92),.clk(clk),.wout(w42_92));
	PE pe42_93(.x(x93),.w(w42_92),.acc(r42_92),.res(r42_93),.clk(clk),.wout(w42_93));
	PE pe42_94(.x(x94),.w(w42_93),.acc(r42_93),.res(r42_94),.clk(clk),.wout(w42_94));
	PE pe42_95(.x(x95),.w(w42_94),.acc(r42_94),.res(r42_95),.clk(clk),.wout(w42_95));
	PE pe42_96(.x(x96),.w(w42_95),.acc(r42_95),.res(r42_96),.clk(clk),.wout(w42_96));
	PE pe42_97(.x(x97),.w(w42_96),.acc(r42_96),.res(r42_97),.clk(clk),.wout(w42_97));
	PE pe42_98(.x(x98),.w(w42_97),.acc(r42_97),.res(r42_98),.clk(clk),.wout(w42_98));
	PE pe42_99(.x(x99),.w(w42_98),.acc(r42_98),.res(r42_99),.clk(clk),.wout(w42_99));
	PE pe42_100(.x(x100),.w(w42_99),.acc(r42_99),.res(r42_100),.clk(clk),.wout(w42_100));
	PE pe42_101(.x(x101),.w(w42_100),.acc(r42_100),.res(r42_101),.clk(clk),.wout(w42_101));
	PE pe42_102(.x(x102),.w(w42_101),.acc(r42_101),.res(r42_102),.clk(clk),.wout(w42_102));
	PE pe42_103(.x(x103),.w(w42_102),.acc(r42_102),.res(r42_103),.clk(clk),.wout(w42_103));
	PE pe42_104(.x(x104),.w(w42_103),.acc(r42_103),.res(r42_104),.clk(clk),.wout(w42_104));
	PE pe42_105(.x(x105),.w(w42_104),.acc(r42_104),.res(r42_105),.clk(clk),.wout(w42_105));
	PE pe42_106(.x(x106),.w(w42_105),.acc(r42_105),.res(r42_106),.clk(clk),.wout(w42_106));
	PE pe42_107(.x(x107),.w(w42_106),.acc(r42_106),.res(r42_107),.clk(clk),.wout(w42_107));
	PE pe42_108(.x(x108),.w(w42_107),.acc(r42_107),.res(r42_108),.clk(clk),.wout(w42_108));
	PE pe42_109(.x(x109),.w(w42_108),.acc(r42_108),.res(r42_109),.clk(clk),.wout(w42_109));
	PE pe42_110(.x(x110),.w(w42_109),.acc(r42_109),.res(r42_110),.clk(clk),.wout(w42_110));
	PE pe42_111(.x(x111),.w(w42_110),.acc(r42_110),.res(r42_111),.clk(clk),.wout(w42_111));
	PE pe42_112(.x(x112),.w(w42_111),.acc(r42_111),.res(r42_112),.clk(clk),.wout(w42_112));
	PE pe42_113(.x(x113),.w(w42_112),.acc(r42_112),.res(r42_113),.clk(clk),.wout(w42_113));
	PE pe42_114(.x(x114),.w(w42_113),.acc(r42_113),.res(r42_114),.clk(clk),.wout(w42_114));
	PE pe42_115(.x(x115),.w(w42_114),.acc(r42_114),.res(r42_115),.clk(clk),.wout(w42_115));
	PE pe42_116(.x(x116),.w(w42_115),.acc(r42_115),.res(r42_116),.clk(clk),.wout(w42_116));
	PE pe42_117(.x(x117),.w(w42_116),.acc(r42_116),.res(r42_117),.clk(clk),.wout(w42_117));
	PE pe42_118(.x(x118),.w(w42_117),.acc(r42_117),.res(r42_118),.clk(clk),.wout(w42_118));
	PE pe42_119(.x(x119),.w(w42_118),.acc(r42_118),.res(r42_119),.clk(clk),.wout(w42_119));
	PE pe42_120(.x(x120),.w(w42_119),.acc(r42_119),.res(r42_120),.clk(clk),.wout(w42_120));
	PE pe42_121(.x(x121),.w(w42_120),.acc(r42_120),.res(r42_121),.clk(clk),.wout(w42_121));
	PE pe42_122(.x(x122),.w(w42_121),.acc(r42_121),.res(r42_122),.clk(clk),.wout(w42_122));
	PE pe42_123(.x(x123),.w(w42_122),.acc(r42_122),.res(r42_123),.clk(clk),.wout(w42_123));
	PE pe42_124(.x(x124),.w(w42_123),.acc(r42_123),.res(r42_124),.clk(clk),.wout(w42_124));
	PE pe42_125(.x(x125),.w(w42_124),.acc(r42_124),.res(r42_125),.clk(clk),.wout(w42_125));
	PE pe42_126(.x(x126),.w(w42_125),.acc(r42_125),.res(r42_126),.clk(clk),.wout(w42_126));
	PE pe42_127(.x(x127),.w(w42_126),.acc(r42_126),.res(result42),.clk(clk),.wout(weight42));

	PE pe43_0(.x(x0),.w(w43),.acc(32'h0),.res(r43_0),.clk(clk),.wout(w43_0));
	PE pe43_1(.x(x1),.w(w43_0),.acc(r43_0),.res(r43_1),.clk(clk),.wout(w43_1));
	PE pe43_2(.x(x2),.w(w43_1),.acc(r43_1),.res(r43_2),.clk(clk),.wout(w43_2));
	PE pe43_3(.x(x3),.w(w43_2),.acc(r43_2),.res(r43_3),.clk(clk),.wout(w43_3));
	PE pe43_4(.x(x4),.w(w43_3),.acc(r43_3),.res(r43_4),.clk(clk),.wout(w43_4));
	PE pe43_5(.x(x5),.w(w43_4),.acc(r43_4),.res(r43_5),.clk(clk),.wout(w43_5));
	PE pe43_6(.x(x6),.w(w43_5),.acc(r43_5),.res(r43_6),.clk(clk),.wout(w43_6));
	PE pe43_7(.x(x7),.w(w43_6),.acc(r43_6),.res(r43_7),.clk(clk),.wout(w43_7));
	PE pe43_8(.x(x8),.w(w43_7),.acc(r43_7),.res(r43_8),.clk(clk),.wout(w43_8));
	PE pe43_9(.x(x9),.w(w43_8),.acc(r43_8),.res(r43_9),.clk(clk),.wout(w43_9));
	PE pe43_10(.x(x10),.w(w43_9),.acc(r43_9),.res(r43_10),.clk(clk),.wout(w43_10));
	PE pe43_11(.x(x11),.w(w43_10),.acc(r43_10),.res(r43_11),.clk(clk),.wout(w43_11));
	PE pe43_12(.x(x12),.w(w43_11),.acc(r43_11),.res(r43_12),.clk(clk),.wout(w43_12));
	PE pe43_13(.x(x13),.w(w43_12),.acc(r43_12),.res(r43_13),.clk(clk),.wout(w43_13));
	PE pe43_14(.x(x14),.w(w43_13),.acc(r43_13),.res(r43_14),.clk(clk),.wout(w43_14));
	PE pe43_15(.x(x15),.w(w43_14),.acc(r43_14),.res(r43_15),.clk(clk),.wout(w43_15));
	PE pe43_16(.x(x16),.w(w43_15),.acc(r43_15),.res(r43_16),.clk(clk),.wout(w43_16));
	PE pe43_17(.x(x17),.w(w43_16),.acc(r43_16),.res(r43_17),.clk(clk),.wout(w43_17));
	PE pe43_18(.x(x18),.w(w43_17),.acc(r43_17),.res(r43_18),.clk(clk),.wout(w43_18));
	PE pe43_19(.x(x19),.w(w43_18),.acc(r43_18),.res(r43_19),.clk(clk),.wout(w43_19));
	PE pe43_20(.x(x20),.w(w43_19),.acc(r43_19),.res(r43_20),.clk(clk),.wout(w43_20));
	PE pe43_21(.x(x21),.w(w43_20),.acc(r43_20),.res(r43_21),.clk(clk),.wout(w43_21));
	PE pe43_22(.x(x22),.w(w43_21),.acc(r43_21),.res(r43_22),.clk(clk),.wout(w43_22));
	PE pe43_23(.x(x23),.w(w43_22),.acc(r43_22),.res(r43_23),.clk(clk),.wout(w43_23));
	PE pe43_24(.x(x24),.w(w43_23),.acc(r43_23),.res(r43_24),.clk(clk),.wout(w43_24));
	PE pe43_25(.x(x25),.w(w43_24),.acc(r43_24),.res(r43_25),.clk(clk),.wout(w43_25));
	PE pe43_26(.x(x26),.w(w43_25),.acc(r43_25),.res(r43_26),.clk(clk),.wout(w43_26));
	PE pe43_27(.x(x27),.w(w43_26),.acc(r43_26),.res(r43_27),.clk(clk),.wout(w43_27));
	PE pe43_28(.x(x28),.w(w43_27),.acc(r43_27),.res(r43_28),.clk(clk),.wout(w43_28));
	PE pe43_29(.x(x29),.w(w43_28),.acc(r43_28),.res(r43_29),.clk(clk),.wout(w43_29));
	PE pe43_30(.x(x30),.w(w43_29),.acc(r43_29),.res(r43_30),.clk(clk),.wout(w43_30));
	PE pe43_31(.x(x31),.w(w43_30),.acc(r43_30),.res(r43_31),.clk(clk),.wout(w43_31));
	PE pe43_32(.x(x32),.w(w43_31),.acc(r43_31),.res(r43_32),.clk(clk),.wout(w43_32));
	PE pe43_33(.x(x33),.w(w43_32),.acc(r43_32),.res(r43_33),.clk(clk),.wout(w43_33));
	PE pe43_34(.x(x34),.w(w43_33),.acc(r43_33),.res(r43_34),.clk(clk),.wout(w43_34));
	PE pe43_35(.x(x35),.w(w43_34),.acc(r43_34),.res(r43_35),.clk(clk),.wout(w43_35));
	PE pe43_36(.x(x36),.w(w43_35),.acc(r43_35),.res(r43_36),.clk(clk),.wout(w43_36));
	PE pe43_37(.x(x37),.w(w43_36),.acc(r43_36),.res(r43_37),.clk(clk),.wout(w43_37));
	PE pe43_38(.x(x38),.w(w43_37),.acc(r43_37),.res(r43_38),.clk(clk),.wout(w43_38));
	PE pe43_39(.x(x39),.w(w43_38),.acc(r43_38),.res(r43_39),.clk(clk),.wout(w43_39));
	PE pe43_40(.x(x40),.w(w43_39),.acc(r43_39),.res(r43_40),.clk(clk),.wout(w43_40));
	PE pe43_41(.x(x41),.w(w43_40),.acc(r43_40),.res(r43_41),.clk(clk),.wout(w43_41));
	PE pe43_42(.x(x42),.w(w43_41),.acc(r43_41),.res(r43_42),.clk(clk),.wout(w43_42));
	PE pe43_43(.x(x43),.w(w43_42),.acc(r43_42),.res(r43_43),.clk(clk),.wout(w43_43));
	PE pe43_44(.x(x44),.w(w43_43),.acc(r43_43),.res(r43_44),.clk(clk),.wout(w43_44));
	PE pe43_45(.x(x45),.w(w43_44),.acc(r43_44),.res(r43_45),.clk(clk),.wout(w43_45));
	PE pe43_46(.x(x46),.w(w43_45),.acc(r43_45),.res(r43_46),.clk(clk),.wout(w43_46));
	PE pe43_47(.x(x47),.w(w43_46),.acc(r43_46),.res(r43_47),.clk(clk),.wout(w43_47));
	PE pe43_48(.x(x48),.w(w43_47),.acc(r43_47),.res(r43_48),.clk(clk),.wout(w43_48));
	PE pe43_49(.x(x49),.w(w43_48),.acc(r43_48),.res(r43_49),.clk(clk),.wout(w43_49));
	PE pe43_50(.x(x50),.w(w43_49),.acc(r43_49),.res(r43_50),.clk(clk),.wout(w43_50));
	PE pe43_51(.x(x51),.w(w43_50),.acc(r43_50),.res(r43_51),.clk(clk),.wout(w43_51));
	PE pe43_52(.x(x52),.w(w43_51),.acc(r43_51),.res(r43_52),.clk(clk),.wout(w43_52));
	PE pe43_53(.x(x53),.w(w43_52),.acc(r43_52),.res(r43_53),.clk(clk),.wout(w43_53));
	PE pe43_54(.x(x54),.w(w43_53),.acc(r43_53),.res(r43_54),.clk(clk),.wout(w43_54));
	PE pe43_55(.x(x55),.w(w43_54),.acc(r43_54),.res(r43_55),.clk(clk),.wout(w43_55));
	PE pe43_56(.x(x56),.w(w43_55),.acc(r43_55),.res(r43_56),.clk(clk),.wout(w43_56));
	PE pe43_57(.x(x57),.w(w43_56),.acc(r43_56),.res(r43_57),.clk(clk),.wout(w43_57));
	PE pe43_58(.x(x58),.w(w43_57),.acc(r43_57),.res(r43_58),.clk(clk),.wout(w43_58));
	PE pe43_59(.x(x59),.w(w43_58),.acc(r43_58),.res(r43_59),.clk(clk),.wout(w43_59));
	PE pe43_60(.x(x60),.w(w43_59),.acc(r43_59),.res(r43_60),.clk(clk),.wout(w43_60));
	PE pe43_61(.x(x61),.w(w43_60),.acc(r43_60),.res(r43_61),.clk(clk),.wout(w43_61));
	PE pe43_62(.x(x62),.w(w43_61),.acc(r43_61),.res(r43_62),.clk(clk),.wout(w43_62));
	PE pe43_63(.x(x63),.w(w43_62),.acc(r43_62),.res(r43_63),.clk(clk),.wout(w43_63));
	PE pe43_64(.x(x64),.w(w43_63),.acc(r43_63),.res(r43_64),.clk(clk),.wout(w43_64));
	PE pe43_65(.x(x65),.w(w43_64),.acc(r43_64),.res(r43_65),.clk(clk),.wout(w43_65));
	PE pe43_66(.x(x66),.w(w43_65),.acc(r43_65),.res(r43_66),.clk(clk),.wout(w43_66));
	PE pe43_67(.x(x67),.w(w43_66),.acc(r43_66),.res(r43_67),.clk(clk),.wout(w43_67));
	PE pe43_68(.x(x68),.w(w43_67),.acc(r43_67),.res(r43_68),.clk(clk),.wout(w43_68));
	PE pe43_69(.x(x69),.w(w43_68),.acc(r43_68),.res(r43_69),.clk(clk),.wout(w43_69));
	PE pe43_70(.x(x70),.w(w43_69),.acc(r43_69),.res(r43_70),.clk(clk),.wout(w43_70));
	PE pe43_71(.x(x71),.w(w43_70),.acc(r43_70),.res(r43_71),.clk(clk),.wout(w43_71));
	PE pe43_72(.x(x72),.w(w43_71),.acc(r43_71),.res(r43_72),.clk(clk),.wout(w43_72));
	PE pe43_73(.x(x73),.w(w43_72),.acc(r43_72),.res(r43_73),.clk(clk),.wout(w43_73));
	PE pe43_74(.x(x74),.w(w43_73),.acc(r43_73),.res(r43_74),.clk(clk),.wout(w43_74));
	PE pe43_75(.x(x75),.w(w43_74),.acc(r43_74),.res(r43_75),.clk(clk),.wout(w43_75));
	PE pe43_76(.x(x76),.w(w43_75),.acc(r43_75),.res(r43_76),.clk(clk),.wout(w43_76));
	PE pe43_77(.x(x77),.w(w43_76),.acc(r43_76),.res(r43_77),.clk(clk),.wout(w43_77));
	PE pe43_78(.x(x78),.w(w43_77),.acc(r43_77),.res(r43_78),.clk(clk),.wout(w43_78));
	PE pe43_79(.x(x79),.w(w43_78),.acc(r43_78),.res(r43_79),.clk(clk),.wout(w43_79));
	PE pe43_80(.x(x80),.w(w43_79),.acc(r43_79),.res(r43_80),.clk(clk),.wout(w43_80));
	PE pe43_81(.x(x81),.w(w43_80),.acc(r43_80),.res(r43_81),.clk(clk),.wout(w43_81));
	PE pe43_82(.x(x82),.w(w43_81),.acc(r43_81),.res(r43_82),.clk(clk),.wout(w43_82));
	PE pe43_83(.x(x83),.w(w43_82),.acc(r43_82),.res(r43_83),.clk(clk),.wout(w43_83));
	PE pe43_84(.x(x84),.w(w43_83),.acc(r43_83),.res(r43_84),.clk(clk),.wout(w43_84));
	PE pe43_85(.x(x85),.w(w43_84),.acc(r43_84),.res(r43_85),.clk(clk),.wout(w43_85));
	PE pe43_86(.x(x86),.w(w43_85),.acc(r43_85),.res(r43_86),.clk(clk),.wout(w43_86));
	PE pe43_87(.x(x87),.w(w43_86),.acc(r43_86),.res(r43_87),.clk(clk),.wout(w43_87));
	PE pe43_88(.x(x88),.w(w43_87),.acc(r43_87),.res(r43_88),.clk(clk),.wout(w43_88));
	PE pe43_89(.x(x89),.w(w43_88),.acc(r43_88),.res(r43_89),.clk(clk),.wout(w43_89));
	PE pe43_90(.x(x90),.w(w43_89),.acc(r43_89),.res(r43_90),.clk(clk),.wout(w43_90));
	PE pe43_91(.x(x91),.w(w43_90),.acc(r43_90),.res(r43_91),.clk(clk),.wout(w43_91));
	PE pe43_92(.x(x92),.w(w43_91),.acc(r43_91),.res(r43_92),.clk(clk),.wout(w43_92));
	PE pe43_93(.x(x93),.w(w43_92),.acc(r43_92),.res(r43_93),.clk(clk),.wout(w43_93));
	PE pe43_94(.x(x94),.w(w43_93),.acc(r43_93),.res(r43_94),.clk(clk),.wout(w43_94));
	PE pe43_95(.x(x95),.w(w43_94),.acc(r43_94),.res(r43_95),.clk(clk),.wout(w43_95));
	PE pe43_96(.x(x96),.w(w43_95),.acc(r43_95),.res(r43_96),.clk(clk),.wout(w43_96));
	PE pe43_97(.x(x97),.w(w43_96),.acc(r43_96),.res(r43_97),.clk(clk),.wout(w43_97));
	PE pe43_98(.x(x98),.w(w43_97),.acc(r43_97),.res(r43_98),.clk(clk),.wout(w43_98));
	PE pe43_99(.x(x99),.w(w43_98),.acc(r43_98),.res(r43_99),.clk(clk),.wout(w43_99));
	PE pe43_100(.x(x100),.w(w43_99),.acc(r43_99),.res(r43_100),.clk(clk),.wout(w43_100));
	PE pe43_101(.x(x101),.w(w43_100),.acc(r43_100),.res(r43_101),.clk(clk),.wout(w43_101));
	PE pe43_102(.x(x102),.w(w43_101),.acc(r43_101),.res(r43_102),.clk(clk),.wout(w43_102));
	PE pe43_103(.x(x103),.w(w43_102),.acc(r43_102),.res(r43_103),.clk(clk),.wout(w43_103));
	PE pe43_104(.x(x104),.w(w43_103),.acc(r43_103),.res(r43_104),.clk(clk),.wout(w43_104));
	PE pe43_105(.x(x105),.w(w43_104),.acc(r43_104),.res(r43_105),.clk(clk),.wout(w43_105));
	PE pe43_106(.x(x106),.w(w43_105),.acc(r43_105),.res(r43_106),.clk(clk),.wout(w43_106));
	PE pe43_107(.x(x107),.w(w43_106),.acc(r43_106),.res(r43_107),.clk(clk),.wout(w43_107));
	PE pe43_108(.x(x108),.w(w43_107),.acc(r43_107),.res(r43_108),.clk(clk),.wout(w43_108));
	PE pe43_109(.x(x109),.w(w43_108),.acc(r43_108),.res(r43_109),.clk(clk),.wout(w43_109));
	PE pe43_110(.x(x110),.w(w43_109),.acc(r43_109),.res(r43_110),.clk(clk),.wout(w43_110));
	PE pe43_111(.x(x111),.w(w43_110),.acc(r43_110),.res(r43_111),.clk(clk),.wout(w43_111));
	PE pe43_112(.x(x112),.w(w43_111),.acc(r43_111),.res(r43_112),.clk(clk),.wout(w43_112));
	PE pe43_113(.x(x113),.w(w43_112),.acc(r43_112),.res(r43_113),.clk(clk),.wout(w43_113));
	PE pe43_114(.x(x114),.w(w43_113),.acc(r43_113),.res(r43_114),.clk(clk),.wout(w43_114));
	PE pe43_115(.x(x115),.w(w43_114),.acc(r43_114),.res(r43_115),.clk(clk),.wout(w43_115));
	PE pe43_116(.x(x116),.w(w43_115),.acc(r43_115),.res(r43_116),.clk(clk),.wout(w43_116));
	PE pe43_117(.x(x117),.w(w43_116),.acc(r43_116),.res(r43_117),.clk(clk),.wout(w43_117));
	PE pe43_118(.x(x118),.w(w43_117),.acc(r43_117),.res(r43_118),.clk(clk),.wout(w43_118));
	PE pe43_119(.x(x119),.w(w43_118),.acc(r43_118),.res(r43_119),.clk(clk),.wout(w43_119));
	PE pe43_120(.x(x120),.w(w43_119),.acc(r43_119),.res(r43_120),.clk(clk),.wout(w43_120));
	PE pe43_121(.x(x121),.w(w43_120),.acc(r43_120),.res(r43_121),.clk(clk),.wout(w43_121));
	PE pe43_122(.x(x122),.w(w43_121),.acc(r43_121),.res(r43_122),.clk(clk),.wout(w43_122));
	PE pe43_123(.x(x123),.w(w43_122),.acc(r43_122),.res(r43_123),.clk(clk),.wout(w43_123));
	PE pe43_124(.x(x124),.w(w43_123),.acc(r43_123),.res(r43_124),.clk(clk),.wout(w43_124));
	PE pe43_125(.x(x125),.w(w43_124),.acc(r43_124),.res(r43_125),.clk(clk),.wout(w43_125));
	PE pe43_126(.x(x126),.w(w43_125),.acc(r43_125),.res(r43_126),.clk(clk),.wout(w43_126));
	PE pe43_127(.x(x127),.w(w43_126),.acc(r43_126),.res(result43),.clk(clk),.wout(weight43));

	PE pe44_0(.x(x0),.w(w44),.acc(32'h0),.res(r44_0),.clk(clk),.wout(w44_0));
	PE pe44_1(.x(x1),.w(w44_0),.acc(r44_0),.res(r44_1),.clk(clk),.wout(w44_1));
	PE pe44_2(.x(x2),.w(w44_1),.acc(r44_1),.res(r44_2),.clk(clk),.wout(w44_2));
	PE pe44_3(.x(x3),.w(w44_2),.acc(r44_2),.res(r44_3),.clk(clk),.wout(w44_3));
	PE pe44_4(.x(x4),.w(w44_3),.acc(r44_3),.res(r44_4),.clk(clk),.wout(w44_4));
	PE pe44_5(.x(x5),.w(w44_4),.acc(r44_4),.res(r44_5),.clk(clk),.wout(w44_5));
	PE pe44_6(.x(x6),.w(w44_5),.acc(r44_5),.res(r44_6),.clk(clk),.wout(w44_6));
	PE pe44_7(.x(x7),.w(w44_6),.acc(r44_6),.res(r44_7),.clk(clk),.wout(w44_7));
	PE pe44_8(.x(x8),.w(w44_7),.acc(r44_7),.res(r44_8),.clk(clk),.wout(w44_8));
	PE pe44_9(.x(x9),.w(w44_8),.acc(r44_8),.res(r44_9),.clk(clk),.wout(w44_9));
	PE pe44_10(.x(x10),.w(w44_9),.acc(r44_9),.res(r44_10),.clk(clk),.wout(w44_10));
	PE pe44_11(.x(x11),.w(w44_10),.acc(r44_10),.res(r44_11),.clk(clk),.wout(w44_11));
	PE pe44_12(.x(x12),.w(w44_11),.acc(r44_11),.res(r44_12),.clk(clk),.wout(w44_12));
	PE pe44_13(.x(x13),.w(w44_12),.acc(r44_12),.res(r44_13),.clk(clk),.wout(w44_13));
	PE pe44_14(.x(x14),.w(w44_13),.acc(r44_13),.res(r44_14),.clk(clk),.wout(w44_14));
	PE pe44_15(.x(x15),.w(w44_14),.acc(r44_14),.res(r44_15),.clk(clk),.wout(w44_15));
	PE pe44_16(.x(x16),.w(w44_15),.acc(r44_15),.res(r44_16),.clk(clk),.wout(w44_16));
	PE pe44_17(.x(x17),.w(w44_16),.acc(r44_16),.res(r44_17),.clk(clk),.wout(w44_17));
	PE pe44_18(.x(x18),.w(w44_17),.acc(r44_17),.res(r44_18),.clk(clk),.wout(w44_18));
	PE pe44_19(.x(x19),.w(w44_18),.acc(r44_18),.res(r44_19),.clk(clk),.wout(w44_19));
	PE pe44_20(.x(x20),.w(w44_19),.acc(r44_19),.res(r44_20),.clk(clk),.wout(w44_20));
	PE pe44_21(.x(x21),.w(w44_20),.acc(r44_20),.res(r44_21),.clk(clk),.wout(w44_21));
	PE pe44_22(.x(x22),.w(w44_21),.acc(r44_21),.res(r44_22),.clk(clk),.wout(w44_22));
	PE pe44_23(.x(x23),.w(w44_22),.acc(r44_22),.res(r44_23),.clk(clk),.wout(w44_23));
	PE pe44_24(.x(x24),.w(w44_23),.acc(r44_23),.res(r44_24),.clk(clk),.wout(w44_24));
	PE pe44_25(.x(x25),.w(w44_24),.acc(r44_24),.res(r44_25),.clk(clk),.wout(w44_25));
	PE pe44_26(.x(x26),.w(w44_25),.acc(r44_25),.res(r44_26),.clk(clk),.wout(w44_26));
	PE pe44_27(.x(x27),.w(w44_26),.acc(r44_26),.res(r44_27),.clk(clk),.wout(w44_27));
	PE pe44_28(.x(x28),.w(w44_27),.acc(r44_27),.res(r44_28),.clk(clk),.wout(w44_28));
	PE pe44_29(.x(x29),.w(w44_28),.acc(r44_28),.res(r44_29),.clk(clk),.wout(w44_29));
	PE pe44_30(.x(x30),.w(w44_29),.acc(r44_29),.res(r44_30),.clk(clk),.wout(w44_30));
	PE pe44_31(.x(x31),.w(w44_30),.acc(r44_30),.res(r44_31),.clk(clk),.wout(w44_31));
	PE pe44_32(.x(x32),.w(w44_31),.acc(r44_31),.res(r44_32),.clk(clk),.wout(w44_32));
	PE pe44_33(.x(x33),.w(w44_32),.acc(r44_32),.res(r44_33),.clk(clk),.wout(w44_33));
	PE pe44_34(.x(x34),.w(w44_33),.acc(r44_33),.res(r44_34),.clk(clk),.wout(w44_34));
	PE pe44_35(.x(x35),.w(w44_34),.acc(r44_34),.res(r44_35),.clk(clk),.wout(w44_35));
	PE pe44_36(.x(x36),.w(w44_35),.acc(r44_35),.res(r44_36),.clk(clk),.wout(w44_36));
	PE pe44_37(.x(x37),.w(w44_36),.acc(r44_36),.res(r44_37),.clk(clk),.wout(w44_37));
	PE pe44_38(.x(x38),.w(w44_37),.acc(r44_37),.res(r44_38),.clk(clk),.wout(w44_38));
	PE pe44_39(.x(x39),.w(w44_38),.acc(r44_38),.res(r44_39),.clk(clk),.wout(w44_39));
	PE pe44_40(.x(x40),.w(w44_39),.acc(r44_39),.res(r44_40),.clk(clk),.wout(w44_40));
	PE pe44_41(.x(x41),.w(w44_40),.acc(r44_40),.res(r44_41),.clk(clk),.wout(w44_41));
	PE pe44_42(.x(x42),.w(w44_41),.acc(r44_41),.res(r44_42),.clk(clk),.wout(w44_42));
	PE pe44_43(.x(x43),.w(w44_42),.acc(r44_42),.res(r44_43),.clk(clk),.wout(w44_43));
	PE pe44_44(.x(x44),.w(w44_43),.acc(r44_43),.res(r44_44),.clk(clk),.wout(w44_44));
	PE pe44_45(.x(x45),.w(w44_44),.acc(r44_44),.res(r44_45),.clk(clk),.wout(w44_45));
	PE pe44_46(.x(x46),.w(w44_45),.acc(r44_45),.res(r44_46),.clk(clk),.wout(w44_46));
	PE pe44_47(.x(x47),.w(w44_46),.acc(r44_46),.res(r44_47),.clk(clk),.wout(w44_47));
	PE pe44_48(.x(x48),.w(w44_47),.acc(r44_47),.res(r44_48),.clk(clk),.wout(w44_48));
	PE pe44_49(.x(x49),.w(w44_48),.acc(r44_48),.res(r44_49),.clk(clk),.wout(w44_49));
	PE pe44_50(.x(x50),.w(w44_49),.acc(r44_49),.res(r44_50),.clk(clk),.wout(w44_50));
	PE pe44_51(.x(x51),.w(w44_50),.acc(r44_50),.res(r44_51),.clk(clk),.wout(w44_51));
	PE pe44_52(.x(x52),.w(w44_51),.acc(r44_51),.res(r44_52),.clk(clk),.wout(w44_52));
	PE pe44_53(.x(x53),.w(w44_52),.acc(r44_52),.res(r44_53),.clk(clk),.wout(w44_53));
	PE pe44_54(.x(x54),.w(w44_53),.acc(r44_53),.res(r44_54),.clk(clk),.wout(w44_54));
	PE pe44_55(.x(x55),.w(w44_54),.acc(r44_54),.res(r44_55),.clk(clk),.wout(w44_55));
	PE pe44_56(.x(x56),.w(w44_55),.acc(r44_55),.res(r44_56),.clk(clk),.wout(w44_56));
	PE pe44_57(.x(x57),.w(w44_56),.acc(r44_56),.res(r44_57),.clk(clk),.wout(w44_57));
	PE pe44_58(.x(x58),.w(w44_57),.acc(r44_57),.res(r44_58),.clk(clk),.wout(w44_58));
	PE pe44_59(.x(x59),.w(w44_58),.acc(r44_58),.res(r44_59),.clk(clk),.wout(w44_59));
	PE pe44_60(.x(x60),.w(w44_59),.acc(r44_59),.res(r44_60),.clk(clk),.wout(w44_60));
	PE pe44_61(.x(x61),.w(w44_60),.acc(r44_60),.res(r44_61),.clk(clk),.wout(w44_61));
	PE pe44_62(.x(x62),.w(w44_61),.acc(r44_61),.res(r44_62),.clk(clk),.wout(w44_62));
	PE pe44_63(.x(x63),.w(w44_62),.acc(r44_62),.res(r44_63),.clk(clk),.wout(w44_63));
	PE pe44_64(.x(x64),.w(w44_63),.acc(r44_63),.res(r44_64),.clk(clk),.wout(w44_64));
	PE pe44_65(.x(x65),.w(w44_64),.acc(r44_64),.res(r44_65),.clk(clk),.wout(w44_65));
	PE pe44_66(.x(x66),.w(w44_65),.acc(r44_65),.res(r44_66),.clk(clk),.wout(w44_66));
	PE pe44_67(.x(x67),.w(w44_66),.acc(r44_66),.res(r44_67),.clk(clk),.wout(w44_67));
	PE pe44_68(.x(x68),.w(w44_67),.acc(r44_67),.res(r44_68),.clk(clk),.wout(w44_68));
	PE pe44_69(.x(x69),.w(w44_68),.acc(r44_68),.res(r44_69),.clk(clk),.wout(w44_69));
	PE pe44_70(.x(x70),.w(w44_69),.acc(r44_69),.res(r44_70),.clk(clk),.wout(w44_70));
	PE pe44_71(.x(x71),.w(w44_70),.acc(r44_70),.res(r44_71),.clk(clk),.wout(w44_71));
	PE pe44_72(.x(x72),.w(w44_71),.acc(r44_71),.res(r44_72),.clk(clk),.wout(w44_72));
	PE pe44_73(.x(x73),.w(w44_72),.acc(r44_72),.res(r44_73),.clk(clk),.wout(w44_73));
	PE pe44_74(.x(x74),.w(w44_73),.acc(r44_73),.res(r44_74),.clk(clk),.wout(w44_74));
	PE pe44_75(.x(x75),.w(w44_74),.acc(r44_74),.res(r44_75),.clk(clk),.wout(w44_75));
	PE pe44_76(.x(x76),.w(w44_75),.acc(r44_75),.res(r44_76),.clk(clk),.wout(w44_76));
	PE pe44_77(.x(x77),.w(w44_76),.acc(r44_76),.res(r44_77),.clk(clk),.wout(w44_77));
	PE pe44_78(.x(x78),.w(w44_77),.acc(r44_77),.res(r44_78),.clk(clk),.wout(w44_78));
	PE pe44_79(.x(x79),.w(w44_78),.acc(r44_78),.res(r44_79),.clk(clk),.wout(w44_79));
	PE pe44_80(.x(x80),.w(w44_79),.acc(r44_79),.res(r44_80),.clk(clk),.wout(w44_80));
	PE pe44_81(.x(x81),.w(w44_80),.acc(r44_80),.res(r44_81),.clk(clk),.wout(w44_81));
	PE pe44_82(.x(x82),.w(w44_81),.acc(r44_81),.res(r44_82),.clk(clk),.wout(w44_82));
	PE pe44_83(.x(x83),.w(w44_82),.acc(r44_82),.res(r44_83),.clk(clk),.wout(w44_83));
	PE pe44_84(.x(x84),.w(w44_83),.acc(r44_83),.res(r44_84),.clk(clk),.wout(w44_84));
	PE pe44_85(.x(x85),.w(w44_84),.acc(r44_84),.res(r44_85),.clk(clk),.wout(w44_85));
	PE pe44_86(.x(x86),.w(w44_85),.acc(r44_85),.res(r44_86),.clk(clk),.wout(w44_86));
	PE pe44_87(.x(x87),.w(w44_86),.acc(r44_86),.res(r44_87),.clk(clk),.wout(w44_87));
	PE pe44_88(.x(x88),.w(w44_87),.acc(r44_87),.res(r44_88),.clk(clk),.wout(w44_88));
	PE pe44_89(.x(x89),.w(w44_88),.acc(r44_88),.res(r44_89),.clk(clk),.wout(w44_89));
	PE pe44_90(.x(x90),.w(w44_89),.acc(r44_89),.res(r44_90),.clk(clk),.wout(w44_90));
	PE pe44_91(.x(x91),.w(w44_90),.acc(r44_90),.res(r44_91),.clk(clk),.wout(w44_91));
	PE pe44_92(.x(x92),.w(w44_91),.acc(r44_91),.res(r44_92),.clk(clk),.wout(w44_92));
	PE pe44_93(.x(x93),.w(w44_92),.acc(r44_92),.res(r44_93),.clk(clk),.wout(w44_93));
	PE pe44_94(.x(x94),.w(w44_93),.acc(r44_93),.res(r44_94),.clk(clk),.wout(w44_94));
	PE pe44_95(.x(x95),.w(w44_94),.acc(r44_94),.res(r44_95),.clk(clk),.wout(w44_95));
	PE pe44_96(.x(x96),.w(w44_95),.acc(r44_95),.res(r44_96),.clk(clk),.wout(w44_96));
	PE pe44_97(.x(x97),.w(w44_96),.acc(r44_96),.res(r44_97),.clk(clk),.wout(w44_97));
	PE pe44_98(.x(x98),.w(w44_97),.acc(r44_97),.res(r44_98),.clk(clk),.wout(w44_98));
	PE pe44_99(.x(x99),.w(w44_98),.acc(r44_98),.res(r44_99),.clk(clk),.wout(w44_99));
	PE pe44_100(.x(x100),.w(w44_99),.acc(r44_99),.res(r44_100),.clk(clk),.wout(w44_100));
	PE pe44_101(.x(x101),.w(w44_100),.acc(r44_100),.res(r44_101),.clk(clk),.wout(w44_101));
	PE pe44_102(.x(x102),.w(w44_101),.acc(r44_101),.res(r44_102),.clk(clk),.wout(w44_102));
	PE pe44_103(.x(x103),.w(w44_102),.acc(r44_102),.res(r44_103),.clk(clk),.wout(w44_103));
	PE pe44_104(.x(x104),.w(w44_103),.acc(r44_103),.res(r44_104),.clk(clk),.wout(w44_104));
	PE pe44_105(.x(x105),.w(w44_104),.acc(r44_104),.res(r44_105),.clk(clk),.wout(w44_105));
	PE pe44_106(.x(x106),.w(w44_105),.acc(r44_105),.res(r44_106),.clk(clk),.wout(w44_106));
	PE pe44_107(.x(x107),.w(w44_106),.acc(r44_106),.res(r44_107),.clk(clk),.wout(w44_107));
	PE pe44_108(.x(x108),.w(w44_107),.acc(r44_107),.res(r44_108),.clk(clk),.wout(w44_108));
	PE pe44_109(.x(x109),.w(w44_108),.acc(r44_108),.res(r44_109),.clk(clk),.wout(w44_109));
	PE pe44_110(.x(x110),.w(w44_109),.acc(r44_109),.res(r44_110),.clk(clk),.wout(w44_110));
	PE pe44_111(.x(x111),.w(w44_110),.acc(r44_110),.res(r44_111),.clk(clk),.wout(w44_111));
	PE pe44_112(.x(x112),.w(w44_111),.acc(r44_111),.res(r44_112),.clk(clk),.wout(w44_112));
	PE pe44_113(.x(x113),.w(w44_112),.acc(r44_112),.res(r44_113),.clk(clk),.wout(w44_113));
	PE pe44_114(.x(x114),.w(w44_113),.acc(r44_113),.res(r44_114),.clk(clk),.wout(w44_114));
	PE pe44_115(.x(x115),.w(w44_114),.acc(r44_114),.res(r44_115),.clk(clk),.wout(w44_115));
	PE pe44_116(.x(x116),.w(w44_115),.acc(r44_115),.res(r44_116),.clk(clk),.wout(w44_116));
	PE pe44_117(.x(x117),.w(w44_116),.acc(r44_116),.res(r44_117),.clk(clk),.wout(w44_117));
	PE pe44_118(.x(x118),.w(w44_117),.acc(r44_117),.res(r44_118),.clk(clk),.wout(w44_118));
	PE pe44_119(.x(x119),.w(w44_118),.acc(r44_118),.res(r44_119),.clk(clk),.wout(w44_119));
	PE pe44_120(.x(x120),.w(w44_119),.acc(r44_119),.res(r44_120),.clk(clk),.wout(w44_120));
	PE pe44_121(.x(x121),.w(w44_120),.acc(r44_120),.res(r44_121),.clk(clk),.wout(w44_121));
	PE pe44_122(.x(x122),.w(w44_121),.acc(r44_121),.res(r44_122),.clk(clk),.wout(w44_122));
	PE pe44_123(.x(x123),.w(w44_122),.acc(r44_122),.res(r44_123),.clk(clk),.wout(w44_123));
	PE pe44_124(.x(x124),.w(w44_123),.acc(r44_123),.res(r44_124),.clk(clk),.wout(w44_124));
	PE pe44_125(.x(x125),.w(w44_124),.acc(r44_124),.res(r44_125),.clk(clk),.wout(w44_125));
	PE pe44_126(.x(x126),.w(w44_125),.acc(r44_125),.res(r44_126),.clk(clk),.wout(w44_126));
	PE pe44_127(.x(x127),.w(w44_126),.acc(r44_126),.res(result44),.clk(clk),.wout(weight44));

	PE pe45_0(.x(x0),.w(w45),.acc(32'h0),.res(r45_0),.clk(clk),.wout(w45_0));
	PE pe45_1(.x(x1),.w(w45_0),.acc(r45_0),.res(r45_1),.clk(clk),.wout(w45_1));
	PE pe45_2(.x(x2),.w(w45_1),.acc(r45_1),.res(r45_2),.clk(clk),.wout(w45_2));
	PE pe45_3(.x(x3),.w(w45_2),.acc(r45_2),.res(r45_3),.clk(clk),.wout(w45_3));
	PE pe45_4(.x(x4),.w(w45_3),.acc(r45_3),.res(r45_4),.clk(clk),.wout(w45_4));
	PE pe45_5(.x(x5),.w(w45_4),.acc(r45_4),.res(r45_5),.clk(clk),.wout(w45_5));
	PE pe45_6(.x(x6),.w(w45_5),.acc(r45_5),.res(r45_6),.clk(clk),.wout(w45_6));
	PE pe45_7(.x(x7),.w(w45_6),.acc(r45_6),.res(r45_7),.clk(clk),.wout(w45_7));
	PE pe45_8(.x(x8),.w(w45_7),.acc(r45_7),.res(r45_8),.clk(clk),.wout(w45_8));
	PE pe45_9(.x(x9),.w(w45_8),.acc(r45_8),.res(r45_9),.clk(clk),.wout(w45_9));
	PE pe45_10(.x(x10),.w(w45_9),.acc(r45_9),.res(r45_10),.clk(clk),.wout(w45_10));
	PE pe45_11(.x(x11),.w(w45_10),.acc(r45_10),.res(r45_11),.clk(clk),.wout(w45_11));
	PE pe45_12(.x(x12),.w(w45_11),.acc(r45_11),.res(r45_12),.clk(clk),.wout(w45_12));
	PE pe45_13(.x(x13),.w(w45_12),.acc(r45_12),.res(r45_13),.clk(clk),.wout(w45_13));
	PE pe45_14(.x(x14),.w(w45_13),.acc(r45_13),.res(r45_14),.clk(clk),.wout(w45_14));
	PE pe45_15(.x(x15),.w(w45_14),.acc(r45_14),.res(r45_15),.clk(clk),.wout(w45_15));
	PE pe45_16(.x(x16),.w(w45_15),.acc(r45_15),.res(r45_16),.clk(clk),.wout(w45_16));
	PE pe45_17(.x(x17),.w(w45_16),.acc(r45_16),.res(r45_17),.clk(clk),.wout(w45_17));
	PE pe45_18(.x(x18),.w(w45_17),.acc(r45_17),.res(r45_18),.clk(clk),.wout(w45_18));
	PE pe45_19(.x(x19),.w(w45_18),.acc(r45_18),.res(r45_19),.clk(clk),.wout(w45_19));
	PE pe45_20(.x(x20),.w(w45_19),.acc(r45_19),.res(r45_20),.clk(clk),.wout(w45_20));
	PE pe45_21(.x(x21),.w(w45_20),.acc(r45_20),.res(r45_21),.clk(clk),.wout(w45_21));
	PE pe45_22(.x(x22),.w(w45_21),.acc(r45_21),.res(r45_22),.clk(clk),.wout(w45_22));
	PE pe45_23(.x(x23),.w(w45_22),.acc(r45_22),.res(r45_23),.clk(clk),.wout(w45_23));
	PE pe45_24(.x(x24),.w(w45_23),.acc(r45_23),.res(r45_24),.clk(clk),.wout(w45_24));
	PE pe45_25(.x(x25),.w(w45_24),.acc(r45_24),.res(r45_25),.clk(clk),.wout(w45_25));
	PE pe45_26(.x(x26),.w(w45_25),.acc(r45_25),.res(r45_26),.clk(clk),.wout(w45_26));
	PE pe45_27(.x(x27),.w(w45_26),.acc(r45_26),.res(r45_27),.clk(clk),.wout(w45_27));
	PE pe45_28(.x(x28),.w(w45_27),.acc(r45_27),.res(r45_28),.clk(clk),.wout(w45_28));
	PE pe45_29(.x(x29),.w(w45_28),.acc(r45_28),.res(r45_29),.clk(clk),.wout(w45_29));
	PE pe45_30(.x(x30),.w(w45_29),.acc(r45_29),.res(r45_30),.clk(clk),.wout(w45_30));
	PE pe45_31(.x(x31),.w(w45_30),.acc(r45_30),.res(r45_31),.clk(clk),.wout(w45_31));
	PE pe45_32(.x(x32),.w(w45_31),.acc(r45_31),.res(r45_32),.clk(clk),.wout(w45_32));
	PE pe45_33(.x(x33),.w(w45_32),.acc(r45_32),.res(r45_33),.clk(clk),.wout(w45_33));
	PE pe45_34(.x(x34),.w(w45_33),.acc(r45_33),.res(r45_34),.clk(clk),.wout(w45_34));
	PE pe45_35(.x(x35),.w(w45_34),.acc(r45_34),.res(r45_35),.clk(clk),.wout(w45_35));
	PE pe45_36(.x(x36),.w(w45_35),.acc(r45_35),.res(r45_36),.clk(clk),.wout(w45_36));
	PE pe45_37(.x(x37),.w(w45_36),.acc(r45_36),.res(r45_37),.clk(clk),.wout(w45_37));
	PE pe45_38(.x(x38),.w(w45_37),.acc(r45_37),.res(r45_38),.clk(clk),.wout(w45_38));
	PE pe45_39(.x(x39),.w(w45_38),.acc(r45_38),.res(r45_39),.clk(clk),.wout(w45_39));
	PE pe45_40(.x(x40),.w(w45_39),.acc(r45_39),.res(r45_40),.clk(clk),.wout(w45_40));
	PE pe45_41(.x(x41),.w(w45_40),.acc(r45_40),.res(r45_41),.clk(clk),.wout(w45_41));
	PE pe45_42(.x(x42),.w(w45_41),.acc(r45_41),.res(r45_42),.clk(clk),.wout(w45_42));
	PE pe45_43(.x(x43),.w(w45_42),.acc(r45_42),.res(r45_43),.clk(clk),.wout(w45_43));
	PE pe45_44(.x(x44),.w(w45_43),.acc(r45_43),.res(r45_44),.clk(clk),.wout(w45_44));
	PE pe45_45(.x(x45),.w(w45_44),.acc(r45_44),.res(r45_45),.clk(clk),.wout(w45_45));
	PE pe45_46(.x(x46),.w(w45_45),.acc(r45_45),.res(r45_46),.clk(clk),.wout(w45_46));
	PE pe45_47(.x(x47),.w(w45_46),.acc(r45_46),.res(r45_47),.clk(clk),.wout(w45_47));
	PE pe45_48(.x(x48),.w(w45_47),.acc(r45_47),.res(r45_48),.clk(clk),.wout(w45_48));
	PE pe45_49(.x(x49),.w(w45_48),.acc(r45_48),.res(r45_49),.clk(clk),.wout(w45_49));
	PE pe45_50(.x(x50),.w(w45_49),.acc(r45_49),.res(r45_50),.clk(clk),.wout(w45_50));
	PE pe45_51(.x(x51),.w(w45_50),.acc(r45_50),.res(r45_51),.clk(clk),.wout(w45_51));
	PE pe45_52(.x(x52),.w(w45_51),.acc(r45_51),.res(r45_52),.clk(clk),.wout(w45_52));
	PE pe45_53(.x(x53),.w(w45_52),.acc(r45_52),.res(r45_53),.clk(clk),.wout(w45_53));
	PE pe45_54(.x(x54),.w(w45_53),.acc(r45_53),.res(r45_54),.clk(clk),.wout(w45_54));
	PE pe45_55(.x(x55),.w(w45_54),.acc(r45_54),.res(r45_55),.clk(clk),.wout(w45_55));
	PE pe45_56(.x(x56),.w(w45_55),.acc(r45_55),.res(r45_56),.clk(clk),.wout(w45_56));
	PE pe45_57(.x(x57),.w(w45_56),.acc(r45_56),.res(r45_57),.clk(clk),.wout(w45_57));
	PE pe45_58(.x(x58),.w(w45_57),.acc(r45_57),.res(r45_58),.clk(clk),.wout(w45_58));
	PE pe45_59(.x(x59),.w(w45_58),.acc(r45_58),.res(r45_59),.clk(clk),.wout(w45_59));
	PE pe45_60(.x(x60),.w(w45_59),.acc(r45_59),.res(r45_60),.clk(clk),.wout(w45_60));
	PE pe45_61(.x(x61),.w(w45_60),.acc(r45_60),.res(r45_61),.clk(clk),.wout(w45_61));
	PE pe45_62(.x(x62),.w(w45_61),.acc(r45_61),.res(r45_62),.clk(clk),.wout(w45_62));
	PE pe45_63(.x(x63),.w(w45_62),.acc(r45_62),.res(r45_63),.clk(clk),.wout(w45_63));
	PE pe45_64(.x(x64),.w(w45_63),.acc(r45_63),.res(r45_64),.clk(clk),.wout(w45_64));
	PE pe45_65(.x(x65),.w(w45_64),.acc(r45_64),.res(r45_65),.clk(clk),.wout(w45_65));
	PE pe45_66(.x(x66),.w(w45_65),.acc(r45_65),.res(r45_66),.clk(clk),.wout(w45_66));
	PE pe45_67(.x(x67),.w(w45_66),.acc(r45_66),.res(r45_67),.clk(clk),.wout(w45_67));
	PE pe45_68(.x(x68),.w(w45_67),.acc(r45_67),.res(r45_68),.clk(clk),.wout(w45_68));
	PE pe45_69(.x(x69),.w(w45_68),.acc(r45_68),.res(r45_69),.clk(clk),.wout(w45_69));
	PE pe45_70(.x(x70),.w(w45_69),.acc(r45_69),.res(r45_70),.clk(clk),.wout(w45_70));
	PE pe45_71(.x(x71),.w(w45_70),.acc(r45_70),.res(r45_71),.clk(clk),.wout(w45_71));
	PE pe45_72(.x(x72),.w(w45_71),.acc(r45_71),.res(r45_72),.clk(clk),.wout(w45_72));
	PE pe45_73(.x(x73),.w(w45_72),.acc(r45_72),.res(r45_73),.clk(clk),.wout(w45_73));
	PE pe45_74(.x(x74),.w(w45_73),.acc(r45_73),.res(r45_74),.clk(clk),.wout(w45_74));
	PE pe45_75(.x(x75),.w(w45_74),.acc(r45_74),.res(r45_75),.clk(clk),.wout(w45_75));
	PE pe45_76(.x(x76),.w(w45_75),.acc(r45_75),.res(r45_76),.clk(clk),.wout(w45_76));
	PE pe45_77(.x(x77),.w(w45_76),.acc(r45_76),.res(r45_77),.clk(clk),.wout(w45_77));
	PE pe45_78(.x(x78),.w(w45_77),.acc(r45_77),.res(r45_78),.clk(clk),.wout(w45_78));
	PE pe45_79(.x(x79),.w(w45_78),.acc(r45_78),.res(r45_79),.clk(clk),.wout(w45_79));
	PE pe45_80(.x(x80),.w(w45_79),.acc(r45_79),.res(r45_80),.clk(clk),.wout(w45_80));
	PE pe45_81(.x(x81),.w(w45_80),.acc(r45_80),.res(r45_81),.clk(clk),.wout(w45_81));
	PE pe45_82(.x(x82),.w(w45_81),.acc(r45_81),.res(r45_82),.clk(clk),.wout(w45_82));
	PE pe45_83(.x(x83),.w(w45_82),.acc(r45_82),.res(r45_83),.clk(clk),.wout(w45_83));
	PE pe45_84(.x(x84),.w(w45_83),.acc(r45_83),.res(r45_84),.clk(clk),.wout(w45_84));
	PE pe45_85(.x(x85),.w(w45_84),.acc(r45_84),.res(r45_85),.clk(clk),.wout(w45_85));
	PE pe45_86(.x(x86),.w(w45_85),.acc(r45_85),.res(r45_86),.clk(clk),.wout(w45_86));
	PE pe45_87(.x(x87),.w(w45_86),.acc(r45_86),.res(r45_87),.clk(clk),.wout(w45_87));
	PE pe45_88(.x(x88),.w(w45_87),.acc(r45_87),.res(r45_88),.clk(clk),.wout(w45_88));
	PE pe45_89(.x(x89),.w(w45_88),.acc(r45_88),.res(r45_89),.clk(clk),.wout(w45_89));
	PE pe45_90(.x(x90),.w(w45_89),.acc(r45_89),.res(r45_90),.clk(clk),.wout(w45_90));
	PE pe45_91(.x(x91),.w(w45_90),.acc(r45_90),.res(r45_91),.clk(clk),.wout(w45_91));
	PE pe45_92(.x(x92),.w(w45_91),.acc(r45_91),.res(r45_92),.clk(clk),.wout(w45_92));
	PE pe45_93(.x(x93),.w(w45_92),.acc(r45_92),.res(r45_93),.clk(clk),.wout(w45_93));
	PE pe45_94(.x(x94),.w(w45_93),.acc(r45_93),.res(r45_94),.clk(clk),.wout(w45_94));
	PE pe45_95(.x(x95),.w(w45_94),.acc(r45_94),.res(r45_95),.clk(clk),.wout(w45_95));
	PE pe45_96(.x(x96),.w(w45_95),.acc(r45_95),.res(r45_96),.clk(clk),.wout(w45_96));
	PE pe45_97(.x(x97),.w(w45_96),.acc(r45_96),.res(r45_97),.clk(clk),.wout(w45_97));
	PE pe45_98(.x(x98),.w(w45_97),.acc(r45_97),.res(r45_98),.clk(clk),.wout(w45_98));
	PE pe45_99(.x(x99),.w(w45_98),.acc(r45_98),.res(r45_99),.clk(clk),.wout(w45_99));
	PE pe45_100(.x(x100),.w(w45_99),.acc(r45_99),.res(r45_100),.clk(clk),.wout(w45_100));
	PE pe45_101(.x(x101),.w(w45_100),.acc(r45_100),.res(r45_101),.clk(clk),.wout(w45_101));
	PE pe45_102(.x(x102),.w(w45_101),.acc(r45_101),.res(r45_102),.clk(clk),.wout(w45_102));
	PE pe45_103(.x(x103),.w(w45_102),.acc(r45_102),.res(r45_103),.clk(clk),.wout(w45_103));
	PE pe45_104(.x(x104),.w(w45_103),.acc(r45_103),.res(r45_104),.clk(clk),.wout(w45_104));
	PE pe45_105(.x(x105),.w(w45_104),.acc(r45_104),.res(r45_105),.clk(clk),.wout(w45_105));
	PE pe45_106(.x(x106),.w(w45_105),.acc(r45_105),.res(r45_106),.clk(clk),.wout(w45_106));
	PE pe45_107(.x(x107),.w(w45_106),.acc(r45_106),.res(r45_107),.clk(clk),.wout(w45_107));
	PE pe45_108(.x(x108),.w(w45_107),.acc(r45_107),.res(r45_108),.clk(clk),.wout(w45_108));
	PE pe45_109(.x(x109),.w(w45_108),.acc(r45_108),.res(r45_109),.clk(clk),.wout(w45_109));
	PE pe45_110(.x(x110),.w(w45_109),.acc(r45_109),.res(r45_110),.clk(clk),.wout(w45_110));
	PE pe45_111(.x(x111),.w(w45_110),.acc(r45_110),.res(r45_111),.clk(clk),.wout(w45_111));
	PE pe45_112(.x(x112),.w(w45_111),.acc(r45_111),.res(r45_112),.clk(clk),.wout(w45_112));
	PE pe45_113(.x(x113),.w(w45_112),.acc(r45_112),.res(r45_113),.clk(clk),.wout(w45_113));
	PE pe45_114(.x(x114),.w(w45_113),.acc(r45_113),.res(r45_114),.clk(clk),.wout(w45_114));
	PE pe45_115(.x(x115),.w(w45_114),.acc(r45_114),.res(r45_115),.clk(clk),.wout(w45_115));
	PE pe45_116(.x(x116),.w(w45_115),.acc(r45_115),.res(r45_116),.clk(clk),.wout(w45_116));
	PE pe45_117(.x(x117),.w(w45_116),.acc(r45_116),.res(r45_117),.clk(clk),.wout(w45_117));
	PE pe45_118(.x(x118),.w(w45_117),.acc(r45_117),.res(r45_118),.clk(clk),.wout(w45_118));
	PE pe45_119(.x(x119),.w(w45_118),.acc(r45_118),.res(r45_119),.clk(clk),.wout(w45_119));
	PE pe45_120(.x(x120),.w(w45_119),.acc(r45_119),.res(r45_120),.clk(clk),.wout(w45_120));
	PE pe45_121(.x(x121),.w(w45_120),.acc(r45_120),.res(r45_121),.clk(clk),.wout(w45_121));
	PE pe45_122(.x(x122),.w(w45_121),.acc(r45_121),.res(r45_122),.clk(clk),.wout(w45_122));
	PE pe45_123(.x(x123),.w(w45_122),.acc(r45_122),.res(r45_123),.clk(clk),.wout(w45_123));
	PE pe45_124(.x(x124),.w(w45_123),.acc(r45_123),.res(r45_124),.clk(clk),.wout(w45_124));
	PE pe45_125(.x(x125),.w(w45_124),.acc(r45_124),.res(r45_125),.clk(clk),.wout(w45_125));
	PE pe45_126(.x(x126),.w(w45_125),.acc(r45_125),.res(r45_126),.clk(clk),.wout(w45_126));
	PE pe45_127(.x(x127),.w(w45_126),.acc(r45_126),.res(result45),.clk(clk),.wout(weight45));

	PE pe46_0(.x(x0),.w(w46),.acc(32'h0),.res(r46_0),.clk(clk),.wout(w46_0));
	PE pe46_1(.x(x1),.w(w46_0),.acc(r46_0),.res(r46_1),.clk(clk),.wout(w46_1));
	PE pe46_2(.x(x2),.w(w46_1),.acc(r46_1),.res(r46_2),.clk(clk),.wout(w46_2));
	PE pe46_3(.x(x3),.w(w46_2),.acc(r46_2),.res(r46_3),.clk(clk),.wout(w46_3));
	PE pe46_4(.x(x4),.w(w46_3),.acc(r46_3),.res(r46_4),.clk(clk),.wout(w46_4));
	PE pe46_5(.x(x5),.w(w46_4),.acc(r46_4),.res(r46_5),.clk(clk),.wout(w46_5));
	PE pe46_6(.x(x6),.w(w46_5),.acc(r46_5),.res(r46_6),.clk(clk),.wout(w46_6));
	PE pe46_7(.x(x7),.w(w46_6),.acc(r46_6),.res(r46_7),.clk(clk),.wout(w46_7));
	PE pe46_8(.x(x8),.w(w46_7),.acc(r46_7),.res(r46_8),.clk(clk),.wout(w46_8));
	PE pe46_9(.x(x9),.w(w46_8),.acc(r46_8),.res(r46_9),.clk(clk),.wout(w46_9));
	PE pe46_10(.x(x10),.w(w46_9),.acc(r46_9),.res(r46_10),.clk(clk),.wout(w46_10));
	PE pe46_11(.x(x11),.w(w46_10),.acc(r46_10),.res(r46_11),.clk(clk),.wout(w46_11));
	PE pe46_12(.x(x12),.w(w46_11),.acc(r46_11),.res(r46_12),.clk(clk),.wout(w46_12));
	PE pe46_13(.x(x13),.w(w46_12),.acc(r46_12),.res(r46_13),.clk(clk),.wout(w46_13));
	PE pe46_14(.x(x14),.w(w46_13),.acc(r46_13),.res(r46_14),.clk(clk),.wout(w46_14));
	PE pe46_15(.x(x15),.w(w46_14),.acc(r46_14),.res(r46_15),.clk(clk),.wout(w46_15));
	PE pe46_16(.x(x16),.w(w46_15),.acc(r46_15),.res(r46_16),.clk(clk),.wout(w46_16));
	PE pe46_17(.x(x17),.w(w46_16),.acc(r46_16),.res(r46_17),.clk(clk),.wout(w46_17));
	PE pe46_18(.x(x18),.w(w46_17),.acc(r46_17),.res(r46_18),.clk(clk),.wout(w46_18));
	PE pe46_19(.x(x19),.w(w46_18),.acc(r46_18),.res(r46_19),.clk(clk),.wout(w46_19));
	PE pe46_20(.x(x20),.w(w46_19),.acc(r46_19),.res(r46_20),.clk(clk),.wout(w46_20));
	PE pe46_21(.x(x21),.w(w46_20),.acc(r46_20),.res(r46_21),.clk(clk),.wout(w46_21));
	PE pe46_22(.x(x22),.w(w46_21),.acc(r46_21),.res(r46_22),.clk(clk),.wout(w46_22));
	PE pe46_23(.x(x23),.w(w46_22),.acc(r46_22),.res(r46_23),.clk(clk),.wout(w46_23));
	PE pe46_24(.x(x24),.w(w46_23),.acc(r46_23),.res(r46_24),.clk(clk),.wout(w46_24));
	PE pe46_25(.x(x25),.w(w46_24),.acc(r46_24),.res(r46_25),.clk(clk),.wout(w46_25));
	PE pe46_26(.x(x26),.w(w46_25),.acc(r46_25),.res(r46_26),.clk(clk),.wout(w46_26));
	PE pe46_27(.x(x27),.w(w46_26),.acc(r46_26),.res(r46_27),.clk(clk),.wout(w46_27));
	PE pe46_28(.x(x28),.w(w46_27),.acc(r46_27),.res(r46_28),.clk(clk),.wout(w46_28));
	PE pe46_29(.x(x29),.w(w46_28),.acc(r46_28),.res(r46_29),.clk(clk),.wout(w46_29));
	PE pe46_30(.x(x30),.w(w46_29),.acc(r46_29),.res(r46_30),.clk(clk),.wout(w46_30));
	PE pe46_31(.x(x31),.w(w46_30),.acc(r46_30),.res(r46_31),.clk(clk),.wout(w46_31));
	PE pe46_32(.x(x32),.w(w46_31),.acc(r46_31),.res(r46_32),.clk(clk),.wout(w46_32));
	PE pe46_33(.x(x33),.w(w46_32),.acc(r46_32),.res(r46_33),.clk(clk),.wout(w46_33));
	PE pe46_34(.x(x34),.w(w46_33),.acc(r46_33),.res(r46_34),.clk(clk),.wout(w46_34));
	PE pe46_35(.x(x35),.w(w46_34),.acc(r46_34),.res(r46_35),.clk(clk),.wout(w46_35));
	PE pe46_36(.x(x36),.w(w46_35),.acc(r46_35),.res(r46_36),.clk(clk),.wout(w46_36));
	PE pe46_37(.x(x37),.w(w46_36),.acc(r46_36),.res(r46_37),.clk(clk),.wout(w46_37));
	PE pe46_38(.x(x38),.w(w46_37),.acc(r46_37),.res(r46_38),.clk(clk),.wout(w46_38));
	PE pe46_39(.x(x39),.w(w46_38),.acc(r46_38),.res(r46_39),.clk(clk),.wout(w46_39));
	PE pe46_40(.x(x40),.w(w46_39),.acc(r46_39),.res(r46_40),.clk(clk),.wout(w46_40));
	PE pe46_41(.x(x41),.w(w46_40),.acc(r46_40),.res(r46_41),.clk(clk),.wout(w46_41));
	PE pe46_42(.x(x42),.w(w46_41),.acc(r46_41),.res(r46_42),.clk(clk),.wout(w46_42));
	PE pe46_43(.x(x43),.w(w46_42),.acc(r46_42),.res(r46_43),.clk(clk),.wout(w46_43));
	PE pe46_44(.x(x44),.w(w46_43),.acc(r46_43),.res(r46_44),.clk(clk),.wout(w46_44));
	PE pe46_45(.x(x45),.w(w46_44),.acc(r46_44),.res(r46_45),.clk(clk),.wout(w46_45));
	PE pe46_46(.x(x46),.w(w46_45),.acc(r46_45),.res(r46_46),.clk(clk),.wout(w46_46));
	PE pe46_47(.x(x47),.w(w46_46),.acc(r46_46),.res(r46_47),.clk(clk),.wout(w46_47));
	PE pe46_48(.x(x48),.w(w46_47),.acc(r46_47),.res(r46_48),.clk(clk),.wout(w46_48));
	PE pe46_49(.x(x49),.w(w46_48),.acc(r46_48),.res(r46_49),.clk(clk),.wout(w46_49));
	PE pe46_50(.x(x50),.w(w46_49),.acc(r46_49),.res(r46_50),.clk(clk),.wout(w46_50));
	PE pe46_51(.x(x51),.w(w46_50),.acc(r46_50),.res(r46_51),.clk(clk),.wout(w46_51));
	PE pe46_52(.x(x52),.w(w46_51),.acc(r46_51),.res(r46_52),.clk(clk),.wout(w46_52));
	PE pe46_53(.x(x53),.w(w46_52),.acc(r46_52),.res(r46_53),.clk(clk),.wout(w46_53));
	PE pe46_54(.x(x54),.w(w46_53),.acc(r46_53),.res(r46_54),.clk(clk),.wout(w46_54));
	PE pe46_55(.x(x55),.w(w46_54),.acc(r46_54),.res(r46_55),.clk(clk),.wout(w46_55));
	PE pe46_56(.x(x56),.w(w46_55),.acc(r46_55),.res(r46_56),.clk(clk),.wout(w46_56));
	PE pe46_57(.x(x57),.w(w46_56),.acc(r46_56),.res(r46_57),.clk(clk),.wout(w46_57));
	PE pe46_58(.x(x58),.w(w46_57),.acc(r46_57),.res(r46_58),.clk(clk),.wout(w46_58));
	PE pe46_59(.x(x59),.w(w46_58),.acc(r46_58),.res(r46_59),.clk(clk),.wout(w46_59));
	PE pe46_60(.x(x60),.w(w46_59),.acc(r46_59),.res(r46_60),.clk(clk),.wout(w46_60));
	PE pe46_61(.x(x61),.w(w46_60),.acc(r46_60),.res(r46_61),.clk(clk),.wout(w46_61));
	PE pe46_62(.x(x62),.w(w46_61),.acc(r46_61),.res(r46_62),.clk(clk),.wout(w46_62));
	PE pe46_63(.x(x63),.w(w46_62),.acc(r46_62),.res(r46_63),.clk(clk),.wout(w46_63));
	PE pe46_64(.x(x64),.w(w46_63),.acc(r46_63),.res(r46_64),.clk(clk),.wout(w46_64));
	PE pe46_65(.x(x65),.w(w46_64),.acc(r46_64),.res(r46_65),.clk(clk),.wout(w46_65));
	PE pe46_66(.x(x66),.w(w46_65),.acc(r46_65),.res(r46_66),.clk(clk),.wout(w46_66));
	PE pe46_67(.x(x67),.w(w46_66),.acc(r46_66),.res(r46_67),.clk(clk),.wout(w46_67));
	PE pe46_68(.x(x68),.w(w46_67),.acc(r46_67),.res(r46_68),.clk(clk),.wout(w46_68));
	PE pe46_69(.x(x69),.w(w46_68),.acc(r46_68),.res(r46_69),.clk(clk),.wout(w46_69));
	PE pe46_70(.x(x70),.w(w46_69),.acc(r46_69),.res(r46_70),.clk(clk),.wout(w46_70));
	PE pe46_71(.x(x71),.w(w46_70),.acc(r46_70),.res(r46_71),.clk(clk),.wout(w46_71));
	PE pe46_72(.x(x72),.w(w46_71),.acc(r46_71),.res(r46_72),.clk(clk),.wout(w46_72));
	PE pe46_73(.x(x73),.w(w46_72),.acc(r46_72),.res(r46_73),.clk(clk),.wout(w46_73));
	PE pe46_74(.x(x74),.w(w46_73),.acc(r46_73),.res(r46_74),.clk(clk),.wout(w46_74));
	PE pe46_75(.x(x75),.w(w46_74),.acc(r46_74),.res(r46_75),.clk(clk),.wout(w46_75));
	PE pe46_76(.x(x76),.w(w46_75),.acc(r46_75),.res(r46_76),.clk(clk),.wout(w46_76));
	PE pe46_77(.x(x77),.w(w46_76),.acc(r46_76),.res(r46_77),.clk(clk),.wout(w46_77));
	PE pe46_78(.x(x78),.w(w46_77),.acc(r46_77),.res(r46_78),.clk(clk),.wout(w46_78));
	PE pe46_79(.x(x79),.w(w46_78),.acc(r46_78),.res(r46_79),.clk(clk),.wout(w46_79));
	PE pe46_80(.x(x80),.w(w46_79),.acc(r46_79),.res(r46_80),.clk(clk),.wout(w46_80));
	PE pe46_81(.x(x81),.w(w46_80),.acc(r46_80),.res(r46_81),.clk(clk),.wout(w46_81));
	PE pe46_82(.x(x82),.w(w46_81),.acc(r46_81),.res(r46_82),.clk(clk),.wout(w46_82));
	PE pe46_83(.x(x83),.w(w46_82),.acc(r46_82),.res(r46_83),.clk(clk),.wout(w46_83));
	PE pe46_84(.x(x84),.w(w46_83),.acc(r46_83),.res(r46_84),.clk(clk),.wout(w46_84));
	PE pe46_85(.x(x85),.w(w46_84),.acc(r46_84),.res(r46_85),.clk(clk),.wout(w46_85));
	PE pe46_86(.x(x86),.w(w46_85),.acc(r46_85),.res(r46_86),.clk(clk),.wout(w46_86));
	PE pe46_87(.x(x87),.w(w46_86),.acc(r46_86),.res(r46_87),.clk(clk),.wout(w46_87));
	PE pe46_88(.x(x88),.w(w46_87),.acc(r46_87),.res(r46_88),.clk(clk),.wout(w46_88));
	PE pe46_89(.x(x89),.w(w46_88),.acc(r46_88),.res(r46_89),.clk(clk),.wout(w46_89));
	PE pe46_90(.x(x90),.w(w46_89),.acc(r46_89),.res(r46_90),.clk(clk),.wout(w46_90));
	PE pe46_91(.x(x91),.w(w46_90),.acc(r46_90),.res(r46_91),.clk(clk),.wout(w46_91));
	PE pe46_92(.x(x92),.w(w46_91),.acc(r46_91),.res(r46_92),.clk(clk),.wout(w46_92));
	PE pe46_93(.x(x93),.w(w46_92),.acc(r46_92),.res(r46_93),.clk(clk),.wout(w46_93));
	PE pe46_94(.x(x94),.w(w46_93),.acc(r46_93),.res(r46_94),.clk(clk),.wout(w46_94));
	PE pe46_95(.x(x95),.w(w46_94),.acc(r46_94),.res(r46_95),.clk(clk),.wout(w46_95));
	PE pe46_96(.x(x96),.w(w46_95),.acc(r46_95),.res(r46_96),.clk(clk),.wout(w46_96));
	PE pe46_97(.x(x97),.w(w46_96),.acc(r46_96),.res(r46_97),.clk(clk),.wout(w46_97));
	PE pe46_98(.x(x98),.w(w46_97),.acc(r46_97),.res(r46_98),.clk(clk),.wout(w46_98));
	PE pe46_99(.x(x99),.w(w46_98),.acc(r46_98),.res(r46_99),.clk(clk),.wout(w46_99));
	PE pe46_100(.x(x100),.w(w46_99),.acc(r46_99),.res(r46_100),.clk(clk),.wout(w46_100));
	PE pe46_101(.x(x101),.w(w46_100),.acc(r46_100),.res(r46_101),.clk(clk),.wout(w46_101));
	PE pe46_102(.x(x102),.w(w46_101),.acc(r46_101),.res(r46_102),.clk(clk),.wout(w46_102));
	PE pe46_103(.x(x103),.w(w46_102),.acc(r46_102),.res(r46_103),.clk(clk),.wout(w46_103));
	PE pe46_104(.x(x104),.w(w46_103),.acc(r46_103),.res(r46_104),.clk(clk),.wout(w46_104));
	PE pe46_105(.x(x105),.w(w46_104),.acc(r46_104),.res(r46_105),.clk(clk),.wout(w46_105));
	PE pe46_106(.x(x106),.w(w46_105),.acc(r46_105),.res(r46_106),.clk(clk),.wout(w46_106));
	PE pe46_107(.x(x107),.w(w46_106),.acc(r46_106),.res(r46_107),.clk(clk),.wout(w46_107));
	PE pe46_108(.x(x108),.w(w46_107),.acc(r46_107),.res(r46_108),.clk(clk),.wout(w46_108));
	PE pe46_109(.x(x109),.w(w46_108),.acc(r46_108),.res(r46_109),.clk(clk),.wout(w46_109));
	PE pe46_110(.x(x110),.w(w46_109),.acc(r46_109),.res(r46_110),.clk(clk),.wout(w46_110));
	PE pe46_111(.x(x111),.w(w46_110),.acc(r46_110),.res(r46_111),.clk(clk),.wout(w46_111));
	PE pe46_112(.x(x112),.w(w46_111),.acc(r46_111),.res(r46_112),.clk(clk),.wout(w46_112));
	PE pe46_113(.x(x113),.w(w46_112),.acc(r46_112),.res(r46_113),.clk(clk),.wout(w46_113));
	PE pe46_114(.x(x114),.w(w46_113),.acc(r46_113),.res(r46_114),.clk(clk),.wout(w46_114));
	PE pe46_115(.x(x115),.w(w46_114),.acc(r46_114),.res(r46_115),.clk(clk),.wout(w46_115));
	PE pe46_116(.x(x116),.w(w46_115),.acc(r46_115),.res(r46_116),.clk(clk),.wout(w46_116));
	PE pe46_117(.x(x117),.w(w46_116),.acc(r46_116),.res(r46_117),.clk(clk),.wout(w46_117));
	PE pe46_118(.x(x118),.w(w46_117),.acc(r46_117),.res(r46_118),.clk(clk),.wout(w46_118));
	PE pe46_119(.x(x119),.w(w46_118),.acc(r46_118),.res(r46_119),.clk(clk),.wout(w46_119));
	PE pe46_120(.x(x120),.w(w46_119),.acc(r46_119),.res(r46_120),.clk(clk),.wout(w46_120));
	PE pe46_121(.x(x121),.w(w46_120),.acc(r46_120),.res(r46_121),.clk(clk),.wout(w46_121));
	PE pe46_122(.x(x122),.w(w46_121),.acc(r46_121),.res(r46_122),.clk(clk),.wout(w46_122));
	PE pe46_123(.x(x123),.w(w46_122),.acc(r46_122),.res(r46_123),.clk(clk),.wout(w46_123));
	PE pe46_124(.x(x124),.w(w46_123),.acc(r46_123),.res(r46_124),.clk(clk),.wout(w46_124));
	PE pe46_125(.x(x125),.w(w46_124),.acc(r46_124),.res(r46_125),.clk(clk),.wout(w46_125));
	PE pe46_126(.x(x126),.w(w46_125),.acc(r46_125),.res(r46_126),.clk(clk),.wout(w46_126));
	PE pe46_127(.x(x127),.w(w46_126),.acc(r46_126),.res(result46),.clk(clk),.wout(weight46));

	PE pe47_0(.x(x0),.w(w47),.acc(32'h0),.res(r47_0),.clk(clk),.wout(w47_0));
	PE pe47_1(.x(x1),.w(w47_0),.acc(r47_0),.res(r47_1),.clk(clk),.wout(w47_1));
	PE pe47_2(.x(x2),.w(w47_1),.acc(r47_1),.res(r47_2),.clk(clk),.wout(w47_2));
	PE pe47_3(.x(x3),.w(w47_2),.acc(r47_2),.res(r47_3),.clk(clk),.wout(w47_3));
	PE pe47_4(.x(x4),.w(w47_3),.acc(r47_3),.res(r47_4),.clk(clk),.wout(w47_4));
	PE pe47_5(.x(x5),.w(w47_4),.acc(r47_4),.res(r47_5),.clk(clk),.wout(w47_5));
	PE pe47_6(.x(x6),.w(w47_5),.acc(r47_5),.res(r47_6),.clk(clk),.wout(w47_6));
	PE pe47_7(.x(x7),.w(w47_6),.acc(r47_6),.res(r47_7),.clk(clk),.wout(w47_7));
	PE pe47_8(.x(x8),.w(w47_7),.acc(r47_7),.res(r47_8),.clk(clk),.wout(w47_8));
	PE pe47_9(.x(x9),.w(w47_8),.acc(r47_8),.res(r47_9),.clk(clk),.wout(w47_9));
	PE pe47_10(.x(x10),.w(w47_9),.acc(r47_9),.res(r47_10),.clk(clk),.wout(w47_10));
	PE pe47_11(.x(x11),.w(w47_10),.acc(r47_10),.res(r47_11),.clk(clk),.wout(w47_11));
	PE pe47_12(.x(x12),.w(w47_11),.acc(r47_11),.res(r47_12),.clk(clk),.wout(w47_12));
	PE pe47_13(.x(x13),.w(w47_12),.acc(r47_12),.res(r47_13),.clk(clk),.wout(w47_13));
	PE pe47_14(.x(x14),.w(w47_13),.acc(r47_13),.res(r47_14),.clk(clk),.wout(w47_14));
	PE pe47_15(.x(x15),.w(w47_14),.acc(r47_14),.res(r47_15),.clk(clk),.wout(w47_15));
	PE pe47_16(.x(x16),.w(w47_15),.acc(r47_15),.res(r47_16),.clk(clk),.wout(w47_16));
	PE pe47_17(.x(x17),.w(w47_16),.acc(r47_16),.res(r47_17),.clk(clk),.wout(w47_17));
	PE pe47_18(.x(x18),.w(w47_17),.acc(r47_17),.res(r47_18),.clk(clk),.wout(w47_18));
	PE pe47_19(.x(x19),.w(w47_18),.acc(r47_18),.res(r47_19),.clk(clk),.wout(w47_19));
	PE pe47_20(.x(x20),.w(w47_19),.acc(r47_19),.res(r47_20),.clk(clk),.wout(w47_20));
	PE pe47_21(.x(x21),.w(w47_20),.acc(r47_20),.res(r47_21),.clk(clk),.wout(w47_21));
	PE pe47_22(.x(x22),.w(w47_21),.acc(r47_21),.res(r47_22),.clk(clk),.wout(w47_22));
	PE pe47_23(.x(x23),.w(w47_22),.acc(r47_22),.res(r47_23),.clk(clk),.wout(w47_23));
	PE pe47_24(.x(x24),.w(w47_23),.acc(r47_23),.res(r47_24),.clk(clk),.wout(w47_24));
	PE pe47_25(.x(x25),.w(w47_24),.acc(r47_24),.res(r47_25),.clk(clk),.wout(w47_25));
	PE pe47_26(.x(x26),.w(w47_25),.acc(r47_25),.res(r47_26),.clk(clk),.wout(w47_26));
	PE pe47_27(.x(x27),.w(w47_26),.acc(r47_26),.res(r47_27),.clk(clk),.wout(w47_27));
	PE pe47_28(.x(x28),.w(w47_27),.acc(r47_27),.res(r47_28),.clk(clk),.wout(w47_28));
	PE pe47_29(.x(x29),.w(w47_28),.acc(r47_28),.res(r47_29),.clk(clk),.wout(w47_29));
	PE pe47_30(.x(x30),.w(w47_29),.acc(r47_29),.res(r47_30),.clk(clk),.wout(w47_30));
	PE pe47_31(.x(x31),.w(w47_30),.acc(r47_30),.res(r47_31),.clk(clk),.wout(w47_31));
	PE pe47_32(.x(x32),.w(w47_31),.acc(r47_31),.res(r47_32),.clk(clk),.wout(w47_32));
	PE pe47_33(.x(x33),.w(w47_32),.acc(r47_32),.res(r47_33),.clk(clk),.wout(w47_33));
	PE pe47_34(.x(x34),.w(w47_33),.acc(r47_33),.res(r47_34),.clk(clk),.wout(w47_34));
	PE pe47_35(.x(x35),.w(w47_34),.acc(r47_34),.res(r47_35),.clk(clk),.wout(w47_35));
	PE pe47_36(.x(x36),.w(w47_35),.acc(r47_35),.res(r47_36),.clk(clk),.wout(w47_36));
	PE pe47_37(.x(x37),.w(w47_36),.acc(r47_36),.res(r47_37),.clk(clk),.wout(w47_37));
	PE pe47_38(.x(x38),.w(w47_37),.acc(r47_37),.res(r47_38),.clk(clk),.wout(w47_38));
	PE pe47_39(.x(x39),.w(w47_38),.acc(r47_38),.res(r47_39),.clk(clk),.wout(w47_39));
	PE pe47_40(.x(x40),.w(w47_39),.acc(r47_39),.res(r47_40),.clk(clk),.wout(w47_40));
	PE pe47_41(.x(x41),.w(w47_40),.acc(r47_40),.res(r47_41),.clk(clk),.wout(w47_41));
	PE pe47_42(.x(x42),.w(w47_41),.acc(r47_41),.res(r47_42),.clk(clk),.wout(w47_42));
	PE pe47_43(.x(x43),.w(w47_42),.acc(r47_42),.res(r47_43),.clk(clk),.wout(w47_43));
	PE pe47_44(.x(x44),.w(w47_43),.acc(r47_43),.res(r47_44),.clk(clk),.wout(w47_44));
	PE pe47_45(.x(x45),.w(w47_44),.acc(r47_44),.res(r47_45),.clk(clk),.wout(w47_45));
	PE pe47_46(.x(x46),.w(w47_45),.acc(r47_45),.res(r47_46),.clk(clk),.wout(w47_46));
	PE pe47_47(.x(x47),.w(w47_46),.acc(r47_46),.res(r47_47),.clk(clk),.wout(w47_47));
	PE pe47_48(.x(x48),.w(w47_47),.acc(r47_47),.res(r47_48),.clk(clk),.wout(w47_48));
	PE pe47_49(.x(x49),.w(w47_48),.acc(r47_48),.res(r47_49),.clk(clk),.wout(w47_49));
	PE pe47_50(.x(x50),.w(w47_49),.acc(r47_49),.res(r47_50),.clk(clk),.wout(w47_50));
	PE pe47_51(.x(x51),.w(w47_50),.acc(r47_50),.res(r47_51),.clk(clk),.wout(w47_51));
	PE pe47_52(.x(x52),.w(w47_51),.acc(r47_51),.res(r47_52),.clk(clk),.wout(w47_52));
	PE pe47_53(.x(x53),.w(w47_52),.acc(r47_52),.res(r47_53),.clk(clk),.wout(w47_53));
	PE pe47_54(.x(x54),.w(w47_53),.acc(r47_53),.res(r47_54),.clk(clk),.wout(w47_54));
	PE pe47_55(.x(x55),.w(w47_54),.acc(r47_54),.res(r47_55),.clk(clk),.wout(w47_55));
	PE pe47_56(.x(x56),.w(w47_55),.acc(r47_55),.res(r47_56),.clk(clk),.wout(w47_56));
	PE pe47_57(.x(x57),.w(w47_56),.acc(r47_56),.res(r47_57),.clk(clk),.wout(w47_57));
	PE pe47_58(.x(x58),.w(w47_57),.acc(r47_57),.res(r47_58),.clk(clk),.wout(w47_58));
	PE pe47_59(.x(x59),.w(w47_58),.acc(r47_58),.res(r47_59),.clk(clk),.wout(w47_59));
	PE pe47_60(.x(x60),.w(w47_59),.acc(r47_59),.res(r47_60),.clk(clk),.wout(w47_60));
	PE pe47_61(.x(x61),.w(w47_60),.acc(r47_60),.res(r47_61),.clk(clk),.wout(w47_61));
	PE pe47_62(.x(x62),.w(w47_61),.acc(r47_61),.res(r47_62),.clk(clk),.wout(w47_62));
	PE pe47_63(.x(x63),.w(w47_62),.acc(r47_62),.res(r47_63),.clk(clk),.wout(w47_63));
	PE pe47_64(.x(x64),.w(w47_63),.acc(r47_63),.res(r47_64),.clk(clk),.wout(w47_64));
	PE pe47_65(.x(x65),.w(w47_64),.acc(r47_64),.res(r47_65),.clk(clk),.wout(w47_65));
	PE pe47_66(.x(x66),.w(w47_65),.acc(r47_65),.res(r47_66),.clk(clk),.wout(w47_66));
	PE pe47_67(.x(x67),.w(w47_66),.acc(r47_66),.res(r47_67),.clk(clk),.wout(w47_67));
	PE pe47_68(.x(x68),.w(w47_67),.acc(r47_67),.res(r47_68),.clk(clk),.wout(w47_68));
	PE pe47_69(.x(x69),.w(w47_68),.acc(r47_68),.res(r47_69),.clk(clk),.wout(w47_69));
	PE pe47_70(.x(x70),.w(w47_69),.acc(r47_69),.res(r47_70),.clk(clk),.wout(w47_70));
	PE pe47_71(.x(x71),.w(w47_70),.acc(r47_70),.res(r47_71),.clk(clk),.wout(w47_71));
	PE pe47_72(.x(x72),.w(w47_71),.acc(r47_71),.res(r47_72),.clk(clk),.wout(w47_72));
	PE pe47_73(.x(x73),.w(w47_72),.acc(r47_72),.res(r47_73),.clk(clk),.wout(w47_73));
	PE pe47_74(.x(x74),.w(w47_73),.acc(r47_73),.res(r47_74),.clk(clk),.wout(w47_74));
	PE pe47_75(.x(x75),.w(w47_74),.acc(r47_74),.res(r47_75),.clk(clk),.wout(w47_75));
	PE pe47_76(.x(x76),.w(w47_75),.acc(r47_75),.res(r47_76),.clk(clk),.wout(w47_76));
	PE pe47_77(.x(x77),.w(w47_76),.acc(r47_76),.res(r47_77),.clk(clk),.wout(w47_77));
	PE pe47_78(.x(x78),.w(w47_77),.acc(r47_77),.res(r47_78),.clk(clk),.wout(w47_78));
	PE pe47_79(.x(x79),.w(w47_78),.acc(r47_78),.res(r47_79),.clk(clk),.wout(w47_79));
	PE pe47_80(.x(x80),.w(w47_79),.acc(r47_79),.res(r47_80),.clk(clk),.wout(w47_80));
	PE pe47_81(.x(x81),.w(w47_80),.acc(r47_80),.res(r47_81),.clk(clk),.wout(w47_81));
	PE pe47_82(.x(x82),.w(w47_81),.acc(r47_81),.res(r47_82),.clk(clk),.wout(w47_82));
	PE pe47_83(.x(x83),.w(w47_82),.acc(r47_82),.res(r47_83),.clk(clk),.wout(w47_83));
	PE pe47_84(.x(x84),.w(w47_83),.acc(r47_83),.res(r47_84),.clk(clk),.wout(w47_84));
	PE pe47_85(.x(x85),.w(w47_84),.acc(r47_84),.res(r47_85),.clk(clk),.wout(w47_85));
	PE pe47_86(.x(x86),.w(w47_85),.acc(r47_85),.res(r47_86),.clk(clk),.wout(w47_86));
	PE pe47_87(.x(x87),.w(w47_86),.acc(r47_86),.res(r47_87),.clk(clk),.wout(w47_87));
	PE pe47_88(.x(x88),.w(w47_87),.acc(r47_87),.res(r47_88),.clk(clk),.wout(w47_88));
	PE pe47_89(.x(x89),.w(w47_88),.acc(r47_88),.res(r47_89),.clk(clk),.wout(w47_89));
	PE pe47_90(.x(x90),.w(w47_89),.acc(r47_89),.res(r47_90),.clk(clk),.wout(w47_90));
	PE pe47_91(.x(x91),.w(w47_90),.acc(r47_90),.res(r47_91),.clk(clk),.wout(w47_91));
	PE pe47_92(.x(x92),.w(w47_91),.acc(r47_91),.res(r47_92),.clk(clk),.wout(w47_92));
	PE pe47_93(.x(x93),.w(w47_92),.acc(r47_92),.res(r47_93),.clk(clk),.wout(w47_93));
	PE pe47_94(.x(x94),.w(w47_93),.acc(r47_93),.res(r47_94),.clk(clk),.wout(w47_94));
	PE pe47_95(.x(x95),.w(w47_94),.acc(r47_94),.res(r47_95),.clk(clk),.wout(w47_95));
	PE pe47_96(.x(x96),.w(w47_95),.acc(r47_95),.res(r47_96),.clk(clk),.wout(w47_96));
	PE pe47_97(.x(x97),.w(w47_96),.acc(r47_96),.res(r47_97),.clk(clk),.wout(w47_97));
	PE pe47_98(.x(x98),.w(w47_97),.acc(r47_97),.res(r47_98),.clk(clk),.wout(w47_98));
	PE pe47_99(.x(x99),.w(w47_98),.acc(r47_98),.res(r47_99),.clk(clk),.wout(w47_99));
	PE pe47_100(.x(x100),.w(w47_99),.acc(r47_99),.res(r47_100),.clk(clk),.wout(w47_100));
	PE pe47_101(.x(x101),.w(w47_100),.acc(r47_100),.res(r47_101),.clk(clk),.wout(w47_101));
	PE pe47_102(.x(x102),.w(w47_101),.acc(r47_101),.res(r47_102),.clk(clk),.wout(w47_102));
	PE pe47_103(.x(x103),.w(w47_102),.acc(r47_102),.res(r47_103),.clk(clk),.wout(w47_103));
	PE pe47_104(.x(x104),.w(w47_103),.acc(r47_103),.res(r47_104),.clk(clk),.wout(w47_104));
	PE pe47_105(.x(x105),.w(w47_104),.acc(r47_104),.res(r47_105),.clk(clk),.wout(w47_105));
	PE pe47_106(.x(x106),.w(w47_105),.acc(r47_105),.res(r47_106),.clk(clk),.wout(w47_106));
	PE pe47_107(.x(x107),.w(w47_106),.acc(r47_106),.res(r47_107),.clk(clk),.wout(w47_107));
	PE pe47_108(.x(x108),.w(w47_107),.acc(r47_107),.res(r47_108),.clk(clk),.wout(w47_108));
	PE pe47_109(.x(x109),.w(w47_108),.acc(r47_108),.res(r47_109),.clk(clk),.wout(w47_109));
	PE pe47_110(.x(x110),.w(w47_109),.acc(r47_109),.res(r47_110),.clk(clk),.wout(w47_110));
	PE pe47_111(.x(x111),.w(w47_110),.acc(r47_110),.res(r47_111),.clk(clk),.wout(w47_111));
	PE pe47_112(.x(x112),.w(w47_111),.acc(r47_111),.res(r47_112),.clk(clk),.wout(w47_112));
	PE pe47_113(.x(x113),.w(w47_112),.acc(r47_112),.res(r47_113),.clk(clk),.wout(w47_113));
	PE pe47_114(.x(x114),.w(w47_113),.acc(r47_113),.res(r47_114),.clk(clk),.wout(w47_114));
	PE pe47_115(.x(x115),.w(w47_114),.acc(r47_114),.res(r47_115),.clk(clk),.wout(w47_115));
	PE pe47_116(.x(x116),.w(w47_115),.acc(r47_115),.res(r47_116),.clk(clk),.wout(w47_116));
	PE pe47_117(.x(x117),.w(w47_116),.acc(r47_116),.res(r47_117),.clk(clk),.wout(w47_117));
	PE pe47_118(.x(x118),.w(w47_117),.acc(r47_117),.res(r47_118),.clk(clk),.wout(w47_118));
	PE pe47_119(.x(x119),.w(w47_118),.acc(r47_118),.res(r47_119),.clk(clk),.wout(w47_119));
	PE pe47_120(.x(x120),.w(w47_119),.acc(r47_119),.res(r47_120),.clk(clk),.wout(w47_120));
	PE pe47_121(.x(x121),.w(w47_120),.acc(r47_120),.res(r47_121),.clk(clk),.wout(w47_121));
	PE pe47_122(.x(x122),.w(w47_121),.acc(r47_121),.res(r47_122),.clk(clk),.wout(w47_122));
	PE pe47_123(.x(x123),.w(w47_122),.acc(r47_122),.res(r47_123),.clk(clk),.wout(w47_123));
	PE pe47_124(.x(x124),.w(w47_123),.acc(r47_123),.res(r47_124),.clk(clk),.wout(w47_124));
	PE pe47_125(.x(x125),.w(w47_124),.acc(r47_124),.res(r47_125),.clk(clk),.wout(w47_125));
	PE pe47_126(.x(x126),.w(w47_125),.acc(r47_125),.res(r47_126),.clk(clk),.wout(w47_126));
	PE pe47_127(.x(x127),.w(w47_126),.acc(r47_126),.res(result47),.clk(clk),.wout(weight47));

	PE pe48_0(.x(x0),.w(w48),.acc(32'h0),.res(r48_0),.clk(clk),.wout(w48_0));
	PE pe48_1(.x(x1),.w(w48_0),.acc(r48_0),.res(r48_1),.clk(clk),.wout(w48_1));
	PE pe48_2(.x(x2),.w(w48_1),.acc(r48_1),.res(r48_2),.clk(clk),.wout(w48_2));
	PE pe48_3(.x(x3),.w(w48_2),.acc(r48_2),.res(r48_3),.clk(clk),.wout(w48_3));
	PE pe48_4(.x(x4),.w(w48_3),.acc(r48_3),.res(r48_4),.clk(clk),.wout(w48_4));
	PE pe48_5(.x(x5),.w(w48_4),.acc(r48_4),.res(r48_5),.clk(clk),.wout(w48_5));
	PE pe48_6(.x(x6),.w(w48_5),.acc(r48_5),.res(r48_6),.clk(clk),.wout(w48_6));
	PE pe48_7(.x(x7),.w(w48_6),.acc(r48_6),.res(r48_7),.clk(clk),.wout(w48_7));
	PE pe48_8(.x(x8),.w(w48_7),.acc(r48_7),.res(r48_8),.clk(clk),.wout(w48_8));
	PE pe48_9(.x(x9),.w(w48_8),.acc(r48_8),.res(r48_9),.clk(clk),.wout(w48_9));
	PE pe48_10(.x(x10),.w(w48_9),.acc(r48_9),.res(r48_10),.clk(clk),.wout(w48_10));
	PE pe48_11(.x(x11),.w(w48_10),.acc(r48_10),.res(r48_11),.clk(clk),.wout(w48_11));
	PE pe48_12(.x(x12),.w(w48_11),.acc(r48_11),.res(r48_12),.clk(clk),.wout(w48_12));
	PE pe48_13(.x(x13),.w(w48_12),.acc(r48_12),.res(r48_13),.clk(clk),.wout(w48_13));
	PE pe48_14(.x(x14),.w(w48_13),.acc(r48_13),.res(r48_14),.clk(clk),.wout(w48_14));
	PE pe48_15(.x(x15),.w(w48_14),.acc(r48_14),.res(r48_15),.clk(clk),.wout(w48_15));
	PE pe48_16(.x(x16),.w(w48_15),.acc(r48_15),.res(r48_16),.clk(clk),.wout(w48_16));
	PE pe48_17(.x(x17),.w(w48_16),.acc(r48_16),.res(r48_17),.clk(clk),.wout(w48_17));
	PE pe48_18(.x(x18),.w(w48_17),.acc(r48_17),.res(r48_18),.clk(clk),.wout(w48_18));
	PE pe48_19(.x(x19),.w(w48_18),.acc(r48_18),.res(r48_19),.clk(clk),.wout(w48_19));
	PE pe48_20(.x(x20),.w(w48_19),.acc(r48_19),.res(r48_20),.clk(clk),.wout(w48_20));
	PE pe48_21(.x(x21),.w(w48_20),.acc(r48_20),.res(r48_21),.clk(clk),.wout(w48_21));
	PE pe48_22(.x(x22),.w(w48_21),.acc(r48_21),.res(r48_22),.clk(clk),.wout(w48_22));
	PE pe48_23(.x(x23),.w(w48_22),.acc(r48_22),.res(r48_23),.clk(clk),.wout(w48_23));
	PE pe48_24(.x(x24),.w(w48_23),.acc(r48_23),.res(r48_24),.clk(clk),.wout(w48_24));
	PE pe48_25(.x(x25),.w(w48_24),.acc(r48_24),.res(r48_25),.clk(clk),.wout(w48_25));
	PE pe48_26(.x(x26),.w(w48_25),.acc(r48_25),.res(r48_26),.clk(clk),.wout(w48_26));
	PE pe48_27(.x(x27),.w(w48_26),.acc(r48_26),.res(r48_27),.clk(clk),.wout(w48_27));
	PE pe48_28(.x(x28),.w(w48_27),.acc(r48_27),.res(r48_28),.clk(clk),.wout(w48_28));
	PE pe48_29(.x(x29),.w(w48_28),.acc(r48_28),.res(r48_29),.clk(clk),.wout(w48_29));
	PE pe48_30(.x(x30),.w(w48_29),.acc(r48_29),.res(r48_30),.clk(clk),.wout(w48_30));
	PE pe48_31(.x(x31),.w(w48_30),.acc(r48_30),.res(r48_31),.clk(clk),.wout(w48_31));
	PE pe48_32(.x(x32),.w(w48_31),.acc(r48_31),.res(r48_32),.clk(clk),.wout(w48_32));
	PE pe48_33(.x(x33),.w(w48_32),.acc(r48_32),.res(r48_33),.clk(clk),.wout(w48_33));
	PE pe48_34(.x(x34),.w(w48_33),.acc(r48_33),.res(r48_34),.clk(clk),.wout(w48_34));
	PE pe48_35(.x(x35),.w(w48_34),.acc(r48_34),.res(r48_35),.clk(clk),.wout(w48_35));
	PE pe48_36(.x(x36),.w(w48_35),.acc(r48_35),.res(r48_36),.clk(clk),.wout(w48_36));
	PE pe48_37(.x(x37),.w(w48_36),.acc(r48_36),.res(r48_37),.clk(clk),.wout(w48_37));
	PE pe48_38(.x(x38),.w(w48_37),.acc(r48_37),.res(r48_38),.clk(clk),.wout(w48_38));
	PE pe48_39(.x(x39),.w(w48_38),.acc(r48_38),.res(r48_39),.clk(clk),.wout(w48_39));
	PE pe48_40(.x(x40),.w(w48_39),.acc(r48_39),.res(r48_40),.clk(clk),.wout(w48_40));
	PE pe48_41(.x(x41),.w(w48_40),.acc(r48_40),.res(r48_41),.clk(clk),.wout(w48_41));
	PE pe48_42(.x(x42),.w(w48_41),.acc(r48_41),.res(r48_42),.clk(clk),.wout(w48_42));
	PE pe48_43(.x(x43),.w(w48_42),.acc(r48_42),.res(r48_43),.clk(clk),.wout(w48_43));
	PE pe48_44(.x(x44),.w(w48_43),.acc(r48_43),.res(r48_44),.clk(clk),.wout(w48_44));
	PE pe48_45(.x(x45),.w(w48_44),.acc(r48_44),.res(r48_45),.clk(clk),.wout(w48_45));
	PE pe48_46(.x(x46),.w(w48_45),.acc(r48_45),.res(r48_46),.clk(clk),.wout(w48_46));
	PE pe48_47(.x(x47),.w(w48_46),.acc(r48_46),.res(r48_47),.clk(clk),.wout(w48_47));
	PE pe48_48(.x(x48),.w(w48_47),.acc(r48_47),.res(r48_48),.clk(clk),.wout(w48_48));
	PE pe48_49(.x(x49),.w(w48_48),.acc(r48_48),.res(r48_49),.clk(clk),.wout(w48_49));
	PE pe48_50(.x(x50),.w(w48_49),.acc(r48_49),.res(r48_50),.clk(clk),.wout(w48_50));
	PE pe48_51(.x(x51),.w(w48_50),.acc(r48_50),.res(r48_51),.clk(clk),.wout(w48_51));
	PE pe48_52(.x(x52),.w(w48_51),.acc(r48_51),.res(r48_52),.clk(clk),.wout(w48_52));
	PE pe48_53(.x(x53),.w(w48_52),.acc(r48_52),.res(r48_53),.clk(clk),.wout(w48_53));
	PE pe48_54(.x(x54),.w(w48_53),.acc(r48_53),.res(r48_54),.clk(clk),.wout(w48_54));
	PE pe48_55(.x(x55),.w(w48_54),.acc(r48_54),.res(r48_55),.clk(clk),.wout(w48_55));
	PE pe48_56(.x(x56),.w(w48_55),.acc(r48_55),.res(r48_56),.clk(clk),.wout(w48_56));
	PE pe48_57(.x(x57),.w(w48_56),.acc(r48_56),.res(r48_57),.clk(clk),.wout(w48_57));
	PE pe48_58(.x(x58),.w(w48_57),.acc(r48_57),.res(r48_58),.clk(clk),.wout(w48_58));
	PE pe48_59(.x(x59),.w(w48_58),.acc(r48_58),.res(r48_59),.clk(clk),.wout(w48_59));
	PE pe48_60(.x(x60),.w(w48_59),.acc(r48_59),.res(r48_60),.clk(clk),.wout(w48_60));
	PE pe48_61(.x(x61),.w(w48_60),.acc(r48_60),.res(r48_61),.clk(clk),.wout(w48_61));
	PE pe48_62(.x(x62),.w(w48_61),.acc(r48_61),.res(r48_62),.clk(clk),.wout(w48_62));
	PE pe48_63(.x(x63),.w(w48_62),.acc(r48_62),.res(r48_63),.clk(clk),.wout(w48_63));
	PE pe48_64(.x(x64),.w(w48_63),.acc(r48_63),.res(r48_64),.clk(clk),.wout(w48_64));
	PE pe48_65(.x(x65),.w(w48_64),.acc(r48_64),.res(r48_65),.clk(clk),.wout(w48_65));
	PE pe48_66(.x(x66),.w(w48_65),.acc(r48_65),.res(r48_66),.clk(clk),.wout(w48_66));
	PE pe48_67(.x(x67),.w(w48_66),.acc(r48_66),.res(r48_67),.clk(clk),.wout(w48_67));
	PE pe48_68(.x(x68),.w(w48_67),.acc(r48_67),.res(r48_68),.clk(clk),.wout(w48_68));
	PE pe48_69(.x(x69),.w(w48_68),.acc(r48_68),.res(r48_69),.clk(clk),.wout(w48_69));
	PE pe48_70(.x(x70),.w(w48_69),.acc(r48_69),.res(r48_70),.clk(clk),.wout(w48_70));
	PE pe48_71(.x(x71),.w(w48_70),.acc(r48_70),.res(r48_71),.clk(clk),.wout(w48_71));
	PE pe48_72(.x(x72),.w(w48_71),.acc(r48_71),.res(r48_72),.clk(clk),.wout(w48_72));
	PE pe48_73(.x(x73),.w(w48_72),.acc(r48_72),.res(r48_73),.clk(clk),.wout(w48_73));
	PE pe48_74(.x(x74),.w(w48_73),.acc(r48_73),.res(r48_74),.clk(clk),.wout(w48_74));
	PE pe48_75(.x(x75),.w(w48_74),.acc(r48_74),.res(r48_75),.clk(clk),.wout(w48_75));
	PE pe48_76(.x(x76),.w(w48_75),.acc(r48_75),.res(r48_76),.clk(clk),.wout(w48_76));
	PE pe48_77(.x(x77),.w(w48_76),.acc(r48_76),.res(r48_77),.clk(clk),.wout(w48_77));
	PE pe48_78(.x(x78),.w(w48_77),.acc(r48_77),.res(r48_78),.clk(clk),.wout(w48_78));
	PE pe48_79(.x(x79),.w(w48_78),.acc(r48_78),.res(r48_79),.clk(clk),.wout(w48_79));
	PE pe48_80(.x(x80),.w(w48_79),.acc(r48_79),.res(r48_80),.clk(clk),.wout(w48_80));
	PE pe48_81(.x(x81),.w(w48_80),.acc(r48_80),.res(r48_81),.clk(clk),.wout(w48_81));
	PE pe48_82(.x(x82),.w(w48_81),.acc(r48_81),.res(r48_82),.clk(clk),.wout(w48_82));
	PE pe48_83(.x(x83),.w(w48_82),.acc(r48_82),.res(r48_83),.clk(clk),.wout(w48_83));
	PE pe48_84(.x(x84),.w(w48_83),.acc(r48_83),.res(r48_84),.clk(clk),.wout(w48_84));
	PE pe48_85(.x(x85),.w(w48_84),.acc(r48_84),.res(r48_85),.clk(clk),.wout(w48_85));
	PE pe48_86(.x(x86),.w(w48_85),.acc(r48_85),.res(r48_86),.clk(clk),.wout(w48_86));
	PE pe48_87(.x(x87),.w(w48_86),.acc(r48_86),.res(r48_87),.clk(clk),.wout(w48_87));
	PE pe48_88(.x(x88),.w(w48_87),.acc(r48_87),.res(r48_88),.clk(clk),.wout(w48_88));
	PE pe48_89(.x(x89),.w(w48_88),.acc(r48_88),.res(r48_89),.clk(clk),.wout(w48_89));
	PE pe48_90(.x(x90),.w(w48_89),.acc(r48_89),.res(r48_90),.clk(clk),.wout(w48_90));
	PE pe48_91(.x(x91),.w(w48_90),.acc(r48_90),.res(r48_91),.clk(clk),.wout(w48_91));
	PE pe48_92(.x(x92),.w(w48_91),.acc(r48_91),.res(r48_92),.clk(clk),.wout(w48_92));
	PE pe48_93(.x(x93),.w(w48_92),.acc(r48_92),.res(r48_93),.clk(clk),.wout(w48_93));
	PE pe48_94(.x(x94),.w(w48_93),.acc(r48_93),.res(r48_94),.clk(clk),.wout(w48_94));
	PE pe48_95(.x(x95),.w(w48_94),.acc(r48_94),.res(r48_95),.clk(clk),.wout(w48_95));
	PE pe48_96(.x(x96),.w(w48_95),.acc(r48_95),.res(r48_96),.clk(clk),.wout(w48_96));
	PE pe48_97(.x(x97),.w(w48_96),.acc(r48_96),.res(r48_97),.clk(clk),.wout(w48_97));
	PE pe48_98(.x(x98),.w(w48_97),.acc(r48_97),.res(r48_98),.clk(clk),.wout(w48_98));
	PE pe48_99(.x(x99),.w(w48_98),.acc(r48_98),.res(r48_99),.clk(clk),.wout(w48_99));
	PE pe48_100(.x(x100),.w(w48_99),.acc(r48_99),.res(r48_100),.clk(clk),.wout(w48_100));
	PE pe48_101(.x(x101),.w(w48_100),.acc(r48_100),.res(r48_101),.clk(clk),.wout(w48_101));
	PE pe48_102(.x(x102),.w(w48_101),.acc(r48_101),.res(r48_102),.clk(clk),.wout(w48_102));
	PE pe48_103(.x(x103),.w(w48_102),.acc(r48_102),.res(r48_103),.clk(clk),.wout(w48_103));
	PE pe48_104(.x(x104),.w(w48_103),.acc(r48_103),.res(r48_104),.clk(clk),.wout(w48_104));
	PE pe48_105(.x(x105),.w(w48_104),.acc(r48_104),.res(r48_105),.clk(clk),.wout(w48_105));
	PE pe48_106(.x(x106),.w(w48_105),.acc(r48_105),.res(r48_106),.clk(clk),.wout(w48_106));
	PE pe48_107(.x(x107),.w(w48_106),.acc(r48_106),.res(r48_107),.clk(clk),.wout(w48_107));
	PE pe48_108(.x(x108),.w(w48_107),.acc(r48_107),.res(r48_108),.clk(clk),.wout(w48_108));
	PE pe48_109(.x(x109),.w(w48_108),.acc(r48_108),.res(r48_109),.clk(clk),.wout(w48_109));
	PE pe48_110(.x(x110),.w(w48_109),.acc(r48_109),.res(r48_110),.clk(clk),.wout(w48_110));
	PE pe48_111(.x(x111),.w(w48_110),.acc(r48_110),.res(r48_111),.clk(clk),.wout(w48_111));
	PE pe48_112(.x(x112),.w(w48_111),.acc(r48_111),.res(r48_112),.clk(clk),.wout(w48_112));
	PE pe48_113(.x(x113),.w(w48_112),.acc(r48_112),.res(r48_113),.clk(clk),.wout(w48_113));
	PE pe48_114(.x(x114),.w(w48_113),.acc(r48_113),.res(r48_114),.clk(clk),.wout(w48_114));
	PE pe48_115(.x(x115),.w(w48_114),.acc(r48_114),.res(r48_115),.clk(clk),.wout(w48_115));
	PE pe48_116(.x(x116),.w(w48_115),.acc(r48_115),.res(r48_116),.clk(clk),.wout(w48_116));
	PE pe48_117(.x(x117),.w(w48_116),.acc(r48_116),.res(r48_117),.clk(clk),.wout(w48_117));
	PE pe48_118(.x(x118),.w(w48_117),.acc(r48_117),.res(r48_118),.clk(clk),.wout(w48_118));
	PE pe48_119(.x(x119),.w(w48_118),.acc(r48_118),.res(r48_119),.clk(clk),.wout(w48_119));
	PE pe48_120(.x(x120),.w(w48_119),.acc(r48_119),.res(r48_120),.clk(clk),.wout(w48_120));
	PE pe48_121(.x(x121),.w(w48_120),.acc(r48_120),.res(r48_121),.clk(clk),.wout(w48_121));
	PE pe48_122(.x(x122),.w(w48_121),.acc(r48_121),.res(r48_122),.clk(clk),.wout(w48_122));
	PE pe48_123(.x(x123),.w(w48_122),.acc(r48_122),.res(r48_123),.clk(clk),.wout(w48_123));
	PE pe48_124(.x(x124),.w(w48_123),.acc(r48_123),.res(r48_124),.clk(clk),.wout(w48_124));
	PE pe48_125(.x(x125),.w(w48_124),.acc(r48_124),.res(r48_125),.clk(clk),.wout(w48_125));
	PE pe48_126(.x(x126),.w(w48_125),.acc(r48_125),.res(r48_126),.clk(clk),.wout(w48_126));
	PE pe48_127(.x(x127),.w(w48_126),.acc(r48_126),.res(result48),.clk(clk),.wout(weight48));

	PE pe49_0(.x(x0),.w(w49),.acc(32'h0),.res(r49_0),.clk(clk),.wout(w49_0));
	PE pe49_1(.x(x1),.w(w49_0),.acc(r49_0),.res(r49_1),.clk(clk),.wout(w49_1));
	PE pe49_2(.x(x2),.w(w49_1),.acc(r49_1),.res(r49_2),.clk(clk),.wout(w49_2));
	PE pe49_3(.x(x3),.w(w49_2),.acc(r49_2),.res(r49_3),.clk(clk),.wout(w49_3));
	PE pe49_4(.x(x4),.w(w49_3),.acc(r49_3),.res(r49_4),.clk(clk),.wout(w49_4));
	PE pe49_5(.x(x5),.w(w49_4),.acc(r49_4),.res(r49_5),.clk(clk),.wout(w49_5));
	PE pe49_6(.x(x6),.w(w49_5),.acc(r49_5),.res(r49_6),.clk(clk),.wout(w49_6));
	PE pe49_7(.x(x7),.w(w49_6),.acc(r49_6),.res(r49_7),.clk(clk),.wout(w49_7));
	PE pe49_8(.x(x8),.w(w49_7),.acc(r49_7),.res(r49_8),.clk(clk),.wout(w49_8));
	PE pe49_9(.x(x9),.w(w49_8),.acc(r49_8),.res(r49_9),.clk(clk),.wout(w49_9));
	PE pe49_10(.x(x10),.w(w49_9),.acc(r49_9),.res(r49_10),.clk(clk),.wout(w49_10));
	PE pe49_11(.x(x11),.w(w49_10),.acc(r49_10),.res(r49_11),.clk(clk),.wout(w49_11));
	PE pe49_12(.x(x12),.w(w49_11),.acc(r49_11),.res(r49_12),.clk(clk),.wout(w49_12));
	PE pe49_13(.x(x13),.w(w49_12),.acc(r49_12),.res(r49_13),.clk(clk),.wout(w49_13));
	PE pe49_14(.x(x14),.w(w49_13),.acc(r49_13),.res(r49_14),.clk(clk),.wout(w49_14));
	PE pe49_15(.x(x15),.w(w49_14),.acc(r49_14),.res(r49_15),.clk(clk),.wout(w49_15));
	PE pe49_16(.x(x16),.w(w49_15),.acc(r49_15),.res(r49_16),.clk(clk),.wout(w49_16));
	PE pe49_17(.x(x17),.w(w49_16),.acc(r49_16),.res(r49_17),.clk(clk),.wout(w49_17));
	PE pe49_18(.x(x18),.w(w49_17),.acc(r49_17),.res(r49_18),.clk(clk),.wout(w49_18));
	PE pe49_19(.x(x19),.w(w49_18),.acc(r49_18),.res(r49_19),.clk(clk),.wout(w49_19));
	PE pe49_20(.x(x20),.w(w49_19),.acc(r49_19),.res(r49_20),.clk(clk),.wout(w49_20));
	PE pe49_21(.x(x21),.w(w49_20),.acc(r49_20),.res(r49_21),.clk(clk),.wout(w49_21));
	PE pe49_22(.x(x22),.w(w49_21),.acc(r49_21),.res(r49_22),.clk(clk),.wout(w49_22));
	PE pe49_23(.x(x23),.w(w49_22),.acc(r49_22),.res(r49_23),.clk(clk),.wout(w49_23));
	PE pe49_24(.x(x24),.w(w49_23),.acc(r49_23),.res(r49_24),.clk(clk),.wout(w49_24));
	PE pe49_25(.x(x25),.w(w49_24),.acc(r49_24),.res(r49_25),.clk(clk),.wout(w49_25));
	PE pe49_26(.x(x26),.w(w49_25),.acc(r49_25),.res(r49_26),.clk(clk),.wout(w49_26));
	PE pe49_27(.x(x27),.w(w49_26),.acc(r49_26),.res(r49_27),.clk(clk),.wout(w49_27));
	PE pe49_28(.x(x28),.w(w49_27),.acc(r49_27),.res(r49_28),.clk(clk),.wout(w49_28));
	PE pe49_29(.x(x29),.w(w49_28),.acc(r49_28),.res(r49_29),.clk(clk),.wout(w49_29));
	PE pe49_30(.x(x30),.w(w49_29),.acc(r49_29),.res(r49_30),.clk(clk),.wout(w49_30));
	PE pe49_31(.x(x31),.w(w49_30),.acc(r49_30),.res(r49_31),.clk(clk),.wout(w49_31));
	PE pe49_32(.x(x32),.w(w49_31),.acc(r49_31),.res(r49_32),.clk(clk),.wout(w49_32));
	PE pe49_33(.x(x33),.w(w49_32),.acc(r49_32),.res(r49_33),.clk(clk),.wout(w49_33));
	PE pe49_34(.x(x34),.w(w49_33),.acc(r49_33),.res(r49_34),.clk(clk),.wout(w49_34));
	PE pe49_35(.x(x35),.w(w49_34),.acc(r49_34),.res(r49_35),.clk(clk),.wout(w49_35));
	PE pe49_36(.x(x36),.w(w49_35),.acc(r49_35),.res(r49_36),.clk(clk),.wout(w49_36));
	PE pe49_37(.x(x37),.w(w49_36),.acc(r49_36),.res(r49_37),.clk(clk),.wout(w49_37));
	PE pe49_38(.x(x38),.w(w49_37),.acc(r49_37),.res(r49_38),.clk(clk),.wout(w49_38));
	PE pe49_39(.x(x39),.w(w49_38),.acc(r49_38),.res(r49_39),.clk(clk),.wout(w49_39));
	PE pe49_40(.x(x40),.w(w49_39),.acc(r49_39),.res(r49_40),.clk(clk),.wout(w49_40));
	PE pe49_41(.x(x41),.w(w49_40),.acc(r49_40),.res(r49_41),.clk(clk),.wout(w49_41));
	PE pe49_42(.x(x42),.w(w49_41),.acc(r49_41),.res(r49_42),.clk(clk),.wout(w49_42));
	PE pe49_43(.x(x43),.w(w49_42),.acc(r49_42),.res(r49_43),.clk(clk),.wout(w49_43));
	PE pe49_44(.x(x44),.w(w49_43),.acc(r49_43),.res(r49_44),.clk(clk),.wout(w49_44));
	PE pe49_45(.x(x45),.w(w49_44),.acc(r49_44),.res(r49_45),.clk(clk),.wout(w49_45));
	PE pe49_46(.x(x46),.w(w49_45),.acc(r49_45),.res(r49_46),.clk(clk),.wout(w49_46));
	PE pe49_47(.x(x47),.w(w49_46),.acc(r49_46),.res(r49_47),.clk(clk),.wout(w49_47));
	PE pe49_48(.x(x48),.w(w49_47),.acc(r49_47),.res(r49_48),.clk(clk),.wout(w49_48));
	PE pe49_49(.x(x49),.w(w49_48),.acc(r49_48),.res(r49_49),.clk(clk),.wout(w49_49));
	PE pe49_50(.x(x50),.w(w49_49),.acc(r49_49),.res(r49_50),.clk(clk),.wout(w49_50));
	PE pe49_51(.x(x51),.w(w49_50),.acc(r49_50),.res(r49_51),.clk(clk),.wout(w49_51));
	PE pe49_52(.x(x52),.w(w49_51),.acc(r49_51),.res(r49_52),.clk(clk),.wout(w49_52));
	PE pe49_53(.x(x53),.w(w49_52),.acc(r49_52),.res(r49_53),.clk(clk),.wout(w49_53));
	PE pe49_54(.x(x54),.w(w49_53),.acc(r49_53),.res(r49_54),.clk(clk),.wout(w49_54));
	PE pe49_55(.x(x55),.w(w49_54),.acc(r49_54),.res(r49_55),.clk(clk),.wout(w49_55));
	PE pe49_56(.x(x56),.w(w49_55),.acc(r49_55),.res(r49_56),.clk(clk),.wout(w49_56));
	PE pe49_57(.x(x57),.w(w49_56),.acc(r49_56),.res(r49_57),.clk(clk),.wout(w49_57));
	PE pe49_58(.x(x58),.w(w49_57),.acc(r49_57),.res(r49_58),.clk(clk),.wout(w49_58));
	PE pe49_59(.x(x59),.w(w49_58),.acc(r49_58),.res(r49_59),.clk(clk),.wout(w49_59));
	PE pe49_60(.x(x60),.w(w49_59),.acc(r49_59),.res(r49_60),.clk(clk),.wout(w49_60));
	PE pe49_61(.x(x61),.w(w49_60),.acc(r49_60),.res(r49_61),.clk(clk),.wout(w49_61));
	PE pe49_62(.x(x62),.w(w49_61),.acc(r49_61),.res(r49_62),.clk(clk),.wout(w49_62));
	PE pe49_63(.x(x63),.w(w49_62),.acc(r49_62),.res(r49_63),.clk(clk),.wout(w49_63));
	PE pe49_64(.x(x64),.w(w49_63),.acc(r49_63),.res(r49_64),.clk(clk),.wout(w49_64));
	PE pe49_65(.x(x65),.w(w49_64),.acc(r49_64),.res(r49_65),.clk(clk),.wout(w49_65));
	PE pe49_66(.x(x66),.w(w49_65),.acc(r49_65),.res(r49_66),.clk(clk),.wout(w49_66));
	PE pe49_67(.x(x67),.w(w49_66),.acc(r49_66),.res(r49_67),.clk(clk),.wout(w49_67));
	PE pe49_68(.x(x68),.w(w49_67),.acc(r49_67),.res(r49_68),.clk(clk),.wout(w49_68));
	PE pe49_69(.x(x69),.w(w49_68),.acc(r49_68),.res(r49_69),.clk(clk),.wout(w49_69));
	PE pe49_70(.x(x70),.w(w49_69),.acc(r49_69),.res(r49_70),.clk(clk),.wout(w49_70));
	PE pe49_71(.x(x71),.w(w49_70),.acc(r49_70),.res(r49_71),.clk(clk),.wout(w49_71));
	PE pe49_72(.x(x72),.w(w49_71),.acc(r49_71),.res(r49_72),.clk(clk),.wout(w49_72));
	PE pe49_73(.x(x73),.w(w49_72),.acc(r49_72),.res(r49_73),.clk(clk),.wout(w49_73));
	PE pe49_74(.x(x74),.w(w49_73),.acc(r49_73),.res(r49_74),.clk(clk),.wout(w49_74));
	PE pe49_75(.x(x75),.w(w49_74),.acc(r49_74),.res(r49_75),.clk(clk),.wout(w49_75));
	PE pe49_76(.x(x76),.w(w49_75),.acc(r49_75),.res(r49_76),.clk(clk),.wout(w49_76));
	PE pe49_77(.x(x77),.w(w49_76),.acc(r49_76),.res(r49_77),.clk(clk),.wout(w49_77));
	PE pe49_78(.x(x78),.w(w49_77),.acc(r49_77),.res(r49_78),.clk(clk),.wout(w49_78));
	PE pe49_79(.x(x79),.w(w49_78),.acc(r49_78),.res(r49_79),.clk(clk),.wout(w49_79));
	PE pe49_80(.x(x80),.w(w49_79),.acc(r49_79),.res(r49_80),.clk(clk),.wout(w49_80));
	PE pe49_81(.x(x81),.w(w49_80),.acc(r49_80),.res(r49_81),.clk(clk),.wout(w49_81));
	PE pe49_82(.x(x82),.w(w49_81),.acc(r49_81),.res(r49_82),.clk(clk),.wout(w49_82));
	PE pe49_83(.x(x83),.w(w49_82),.acc(r49_82),.res(r49_83),.clk(clk),.wout(w49_83));
	PE pe49_84(.x(x84),.w(w49_83),.acc(r49_83),.res(r49_84),.clk(clk),.wout(w49_84));
	PE pe49_85(.x(x85),.w(w49_84),.acc(r49_84),.res(r49_85),.clk(clk),.wout(w49_85));
	PE pe49_86(.x(x86),.w(w49_85),.acc(r49_85),.res(r49_86),.clk(clk),.wout(w49_86));
	PE pe49_87(.x(x87),.w(w49_86),.acc(r49_86),.res(r49_87),.clk(clk),.wout(w49_87));
	PE pe49_88(.x(x88),.w(w49_87),.acc(r49_87),.res(r49_88),.clk(clk),.wout(w49_88));
	PE pe49_89(.x(x89),.w(w49_88),.acc(r49_88),.res(r49_89),.clk(clk),.wout(w49_89));
	PE pe49_90(.x(x90),.w(w49_89),.acc(r49_89),.res(r49_90),.clk(clk),.wout(w49_90));
	PE pe49_91(.x(x91),.w(w49_90),.acc(r49_90),.res(r49_91),.clk(clk),.wout(w49_91));
	PE pe49_92(.x(x92),.w(w49_91),.acc(r49_91),.res(r49_92),.clk(clk),.wout(w49_92));
	PE pe49_93(.x(x93),.w(w49_92),.acc(r49_92),.res(r49_93),.clk(clk),.wout(w49_93));
	PE pe49_94(.x(x94),.w(w49_93),.acc(r49_93),.res(r49_94),.clk(clk),.wout(w49_94));
	PE pe49_95(.x(x95),.w(w49_94),.acc(r49_94),.res(r49_95),.clk(clk),.wout(w49_95));
	PE pe49_96(.x(x96),.w(w49_95),.acc(r49_95),.res(r49_96),.clk(clk),.wout(w49_96));
	PE pe49_97(.x(x97),.w(w49_96),.acc(r49_96),.res(r49_97),.clk(clk),.wout(w49_97));
	PE pe49_98(.x(x98),.w(w49_97),.acc(r49_97),.res(r49_98),.clk(clk),.wout(w49_98));
	PE pe49_99(.x(x99),.w(w49_98),.acc(r49_98),.res(r49_99),.clk(clk),.wout(w49_99));
	PE pe49_100(.x(x100),.w(w49_99),.acc(r49_99),.res(r49_100),.clk(clk),.wout(w49_100));
	PE pe49_101(.x(x101),.w(w49_100),.acc(r49_100),.res(r49_101),.clk(clk),.wout(w49_101));
	PE pe49_102(.x(x102),.w(w49_101),.acc(r49_101),.res(r49_102),.clk(clk),.wout(w49_102));
	PE pe49_103(.x(x103),.w(w49_102),.acc(r49_102),.res(r49_103),.clk(clk),.wout(w49_103));
	PE pe49_104(.x(x104),.w(w49_103),.acc(r49_103),.res(r49_104),.clk(clk),.wout(w49_104));
	PE pe49_105(.x(x105),.w(w49_104),.acc(r49_104),.res(r49_105),.clk(clk),.wout(w49_105));
	PE pe49_106(.x(x106),.w(w49_105),.acc(r49_105),.res(r49_106),.clk(clk),.wout(w49_106));
	PE pe49_107(.x(x107),.w(w49_106),.acc(r49_106),.res(r49_107),.clk(clk),.wout(w49_107));
	PE pe49_108(.x(x108),.w(w49_107),.acc(r49_107),.res(r49_108),.clk(clk),.wout(w49_108));
	PE pe49_109(.x(x109),.w(w49_108),.acc(r49_108),.res(r49_109),.clk(clk),.wout(w49_109));
	PE pe49_110(.x(x110),.w(w49_109),.acc(r49_109),.res(r49_110),.clk(clk),.wout(w49_110));
	PE pe49_111(.x(x111),.w(w49_110),.acc(r49_110),.res(r49_111),.clk(clk),.wout(w49_111));
	PE pe49_112(.x(x112),.w(w49_111),.acc(r49_111),.res(r49_112),.clk(clk),.wout(w49_112));
	PE pe49_113(.x(x113),.w(w49_112),.acc(r49_112),.res(r49_113),.clk(clk),.wout(w49_113));
	PE pe49_114(.x(x114),.w(w49_113),.acc(r49_113),.res(r49_114),.clk(clk),.wout(w49_114));
	PE pe49_115(.x(x115),.w(w49_114),.acc(r49_114),.res(r49_115),.clk(clk),.wout(w49_115));
	PE pe49_116(.x(x116),.w(w49_115),.acc(r49_115),.res(r49_116),.clk(clk),.wout(w49_116));
	PE pe49_117(.x(x117),.w(w49_116),.acc(r49_116),.res(r49_117),.clk(clk),.wout(w49_117));
	PE pe49_118(.x(x118),.w(w49_117),.acc(r49_117),.res(r49_118),.clk(clk),.wout(w49_118));
	PE pe49_119(.x(x119),.w(w49_118),.acc(r49_118),.res(r49_119),.clk(clk),.wout(w49_119));
	PE pe49_120(.x(x120),.w(w49_119),.acc(r49_119),.res(r49_120),.clk(clk),.wout(w49_120));
	PE pe49_121(.x(x121),.w(w49_120),.acc(r49_120),.res(r49_121),.clk(clk),.wout(w49_121));
	PE pe49_122(.x(x122),.w(w49_121),.acc(r49_121),.res(r49_122),.clk(clk),.wout(w49_122));
	PE pe49_123(.x(x123),.w(w49_122),.acc(r49_122),.res(r49_123),.clk(clk),.wout(w49_123));
	PE pe49_124(.x(x124),.w(w49_123),.acc(r49_123),.res(r49_124),.clk(clk),.wout(w49_124));
	PE pe49_125(.x(x125),.w(w49_124),.acc(r49_124),.res(r49_125),.clk(clk),.wout(w49_125));
	PE pe49_126(.x(x126),.w(w49_125),.acc(r49_125),.res(r49_126),.clk(clk),.wout(w49_126));
	PE pe49_127(.x(x127),.w(w49_126),.acc(r49_126),.res(result49),.clk(clk),.wout(weight49));

	PE pe50_0(.x(x0),.w(w50),.acc(32'h0),.res(r50_0),.clk(clk),.wout(w50_0));
	PE pe50_1(.x(x1),.w(w50_0),.acc(r50_0),.res(r50_1),.clk(clk),.wout(w50_1));
	PE pe50_2(.x(x2),.w(w50_1),.acc(r50_1),.res(r50_2),.clk(clk),.wout(w50_2));
	PE pe50_3(.x(x3),.w(w50_2),.acc(r50_2),.res(r50_3),.clk(clk),.wout(w50_3));
	PE pe50_4(.x(x4),.w(w50_3),.acc(r50_3),.res(r50_4),.clk(clk),.wout(w50_4));
	PE pe50_5(.x(x5),.w(w50_4),.acc(r50_4),.res(r50_5),.clk(clk),.wout(w50_5));
	PE pe50_6(.x(x6),.w(w50_5),.acc(r50_5),.res(r50_6),.clk(clk),.wout(w50_6));
	PE pe50_7(.x(x7),.w(w50_6),.acc(r50_6),.res(r50_7),.clk(clk),.wout(w50_7));
	PE pe50_8(.x(x8),.w(w50_7),.acc(r50_7),.res(r50_8),.clk(clk),.wout(w50_8));
	PE pe50_9(.x(x9),.w(w50_8),.acc(r50_8),.res(r50_9),.clk(clk),.wout(w50_9));
	PE pe50_10(.x(x10),.w(w50_9),.acc(r50_9),.res(r50_10),.clk(clk),.wout(w50_10));
	PE pe50_11(.x(x11),.w(w50_10),.acc(r50_10),.res(r50_11),.clk(clk),.wout(w50_11));
	PE pe50_12(.x(x12),.w(w50_11),.acc(r50_11),.res(r50_12),.clk(clk),.wout(w50_12));
	PE pe50_13(.x(x13),.w(w50_12),.acc(r50_12),.res(r50_13),.clk(clk),.wout(w50_13));
	PE pe50_14(.x(x14),.w(w50_13),.acc(r50_13),.res(r50_14),.clk(clk),.wout(w50_14));
	PE pe50_15(.x(x15),.w(w50_14),.acc(r50_14),.res(r50_15),.clk(clk),.wout(w50_15));
	PE pe50_16(.x(x16),.w(w50_15),.acc(r50_15),.res(r50_16),.clk(clk),.wout(w50_16));
	PE pe50_17(.x(x17),.w(w50_16),.acc(r50_16),.res(r50_17),.clk(clk),.wout(w50_17));
	PE pe50_18(.x(x18),.w(w50_17),.acc(r50_17),.res(r50_18),.clk(clk),.wout(w50_18));
	PE pe50_19(.x(x19),.w(w50_18),.acc(r50_18),.res(r50_19),.clk(clk),.wout(w50_19));
	PE pe50_20(.x(x20),.w(w50_19),.acc(r50_19),.res(r50_20),.clk(clk),.wout(w50_20));
	PE pe50_21(.x(x21),.w(w50_20),.acc(r50_20),.res(r50_21),.clk(clk),.wout(w50_21));
	PE pe50_22(.x(x22),.w(w50_21),.acc(r50_21),.res(r50_22),.clk(clk),.wout(w50_22));
	PE pe50_23(.x(x23),.w(w50_22),.acc(r50_22),.res(r50_23),.clk(clk),.wout(w50_23));
	PE pe50_24(.x(x24),.w(w50_23),.acc(r50_23),.res(r50_24),.clk(clk),.wout(w50_24));
	PE pe50_25(.x(x25),.w(w50_24),.acc(r50_24),.res(r50_25),.clk(clk),.wout(w50_25));
	PE pe50_26(.x(x26),.w(w50_25),.acc(r50_25),.res(r50_26),.clk(clk),.wout(w50_26));
	PE pe50_27(.x(x27),.w(w50_26),.acc(r50_26),.res(r50_27),.clk(clk),.wout(w50_27));
	PE pe50_28(.x(x28),.w(w50_27),.acc(r50_27),.res(r50_28),.clk(clk),.wout(w50_28));
	PE pe50_29(.x(x29),.w(w50_28),.acc(r50_28),.res(r50_29),.clk(clk),.wout(w50_29));
	PE pe50_30(.x(x30),.w(w50_29),.acc(r50_29),.res(r50_30),.clk(clk),.wout(w50_30));
	PE pe50_31(.x(x31),.w(w50_30),.acc(r50_30),.res(r50_31),.clk(clk),.wout(w50_31));
	PE pe50_32(.x(x32),.w(w50_31),.acc(r50_31),.res(r50_32),.clk(clk),.wout(w50_32));
	PE pe50_33(.x(x33),.w(w50_32),.acc(r50_32),.res(r50_33),.clk(clk),.wout(w50_33));
	PE pe50_34(.x(x34),.w(w50_33),.acc(r50_33),.res(r50_34),.clk(clk),.wout(w50_34));
	PE pe50_35(.x(x35),.w(w50_34),.acc(r50_34),.res(r50_35),.clk(clk),.wout(w50_35));
	PE pe50_36(.x(x36),.w(w50_35),.acc(r50_35),.res(r50_36),.clk(clk),.wout(w50_36));
	PE pe50_37(.x(x37),.w(w50_36),.acc(r50_36),.res(r50_37),.clk(clk),.wout(w50_37));
	PE pe50_38(.x(x38),.w(w50_37),.acc(r50_37),.res(r50_38),.clk(clk),.wout(w50_38));
	PE pe50_39(.x(x39),.w(w50_38),.acc(r50_38),.res(r50_39),.clk(clk),.wout(w50_39));
	PE pe50_40(.x(x40),.w(w50_39),.acc(r50_39),.res(r50_40),.clk(clk),.wout(w50_40));
	PE pe50_41(.x(x41),.w(w50_40),.acc(r50_40),.res(r50_41),.clk(clk),.wout(w50_41));
	PE pe50_42(.x(x42),.w(w50_41),.acc(r50_41),.res(r50_42),.clk(clk),.wout(w50_42));
	PE pe50_43(.x(x43),.w(w50_42),.acc(r50_42),.res(r50_43),.clk(clk),.wout(w50_43));
	PE pe50_44(.x(x44),.w(w50_43),.acc(r50_43),.res(r50_44),.clk(clk),.wout(w50_44));
	PE pe50_45(.x(x45),.w(w50_44),.acc(r50_44),.res(r50_45),.clk(clk),.wout(w50_45));
	PE pe50_46(.x(x46),.w(w50_45),.acc(r50_45),.res(r50_46),.clk(clk),.wout(w50_46));
	PE pe50_47(.x(x47),.w(w50_46),.acc(r50_46),.res(r50_47),.clk(clk),.wout(w50_47));
	PE pe50_48(.x(x48),.w(w50_47),.acc(r50_47),.res(r50_48),.clk(clk),.wout(w50_48));
	PE pe50_49(.x(x49),.w(w50_48),.acc(r50_48),.res(r50_49),.clk(clk),.wout(w50_49));
	PE pe50_50(.x(x50),.w(w50_49),.acc(r50_49),.res(r50_50),.clk(clk),.wout(w50_50));
	PE pe50_51(.x(x51),.w(w50_50),.acc(r50_50),.res(r50_51),.clk(clk),.wout(w50_51));
	PE pe50_52(.x(x52),.w(w50_51),.acc(r50_51),.res(r50_52),.clk(clk),.wout(w50_52));
	PE pe50_53(.x(x53),.w(w50_52),.acc(r50_52),.res(r50_53),.clk(clk),.wout(w50_53));
	PE pe50_54(.x(x54),.w(w50_53),.acc(r50_53),.res(r50_54),.clk(clk),.wout(w50_54));
	PE pe50_55(.x(x55),.w(w50_54),.acc(r50_54),.res(r50_55),.clk(clk),.wout(w50_55));
	PE pe50_56(.x(x56),.w(w50_55),.acc(r50_55),.res(r50_56),.clk(clk),.wout(w50_56));
	PE pe50_57(.x(x57),.w(w50_56),.acc(r50_56),.res(r50_57),.clk(clk),.wout(w50_57));
	PE pe50_58(.x(x58),.w(w50_57),.acc(r50_57),.res(r50_58),.clk(clk),.wout(w50_58));
	PE pe50_59(.x(x59),.w(w50_58),.acc(r50_58),.res(r50_59),.clk(clk),.wout(w50_59));
	PE pe50_60(.x(x60),.w(w50_59),.acc(r50_59),.res(r50_60),.clk(clk),.wout(w50_60));
	PE pe50_61(.x(x61),.w(w50_60),.acc(r50_60),.res(r50_61),.clk(clk),.wout(w50_61));
	PE pe50_62(.x(x62),.w(w50_61),.acc(r50_61),.res(r50_62),.clk(clk),.wout(w50_62));
	PE pe50_63(.x(x63),.w(w50_62),.acc(r50_62),.res(r50_63),.clk(clk),.wout(w50_63));
	PE pe50_64(.x(x64),.w(w50_63),.acc(r50_63),.res(r50_64),.clk(clk),.wout(w50_64));
	PE pe50_65(.x(x65),.w(w50_64),.acc(r50_64),.res(r50_65),.clk(clk),.wout(w50_65));
	PE pe50_66(.x(x66),.w(w50_65),.acc(r50_65),.res(r50_66),.clk(clk),.wout(w50_66));
	PE pe50_67(.x(x67),.w(w50_66),.acc(r50_66),.res(r50_67),.clk(clk),.wout(w50_67));
	PE pe50_68(.x(x68),.w(w50_67),.acc(r50_67),.res(r50_68),.clk(clk),.wout(w50_68));
	PE pe50_69(.x(x69),.w(w50_68),.acc(r50_68),.res(r50_69),.clk(clk),.wout(w50_69));
	PE pe50_70(.x(x70),.w(w50_69),.acc(r50_69),.res(r50_70),.clk(clk),.wout(w50_70));
	PE pe50_71(.x(x71),.w(w50_70),.acc(r50_70),.res(r50_71),.clk(clk),.wout(w50_71));
	PE pe50_72(.x(x72),.w(w50_71),.acc(r50_71),.res(r50_72),.clk(clk),.wout(w50_72));
	PE pe50_73(.x(x73),.w(w50_72),.acc(r50_72),.res(r50_73),.clk(clk),.wout(w50_73));
	PE pe50_74(.x(x74),.w(w50_73),.acc(r50_73),.res(r50_74),.clk(clk),.wout(w50_74));
	PE pe50_75(.x(x75),.w(w50_74),.acc(r50_74),.res(r50_75),.clk(clk),.wout(w50_75));
	PE pe50_76(.x(x76),.w(w50_75),.acc(r50_75),.res(r50_76),.clk(clk),.wout(w50_76));
	PE pe50_77(.x(x77),.w(w50_76),.acc(r50_76),.res(r50_77),.clk(clk),.wout(w50_77));
	PE pe50_78(.x(x78),.w(w50_77),.acc(r50_77),.res(r50_78),.clk(clk),.wout(w50_78));
	PE pe50_79(.x(x79),.w(w50_78),.acc(r50_78),.res(r50_79),.clk(clk),.wout(w50_79));
	PE pe50_80(.x(x80),.w(w50_79),.acc(r50_79),.res(r50_80),.clk(clk),.wout(w50_80));
	PE pe50_81(.x(x81),.w(w50_80),.acc(r50_80),.res(r50_81),.clk(clk),.wout(w50_81));
	PE pe50_82(.x(x82),.w(w50_81),.acc(r50_81),.res(r50_82),.clk(clk),.wout(w50_82));
	PE pe50_83(.x(x83),.w(w50_82),.acc(r50_82),.res(r50_83),.clk(clk),.wout(w50_83));
	PE pe50_84(.x(x84),.w(w50_83),.acc(r50_83),.res(r50_84),.clk(clk),.wout(w50_84));
	PE pe50_85(.x(x85),.w(w50_84),.acc(r50_84),.res(r50_85),.clk(clk),.wout(w50_85));
	PE pe50_86(.x(x86),.w(w50_85),.acc(r50_85),.res(r50_86),.clk(clk),.wout(w50_86));
	PE pe50_87(.x(x87),.w(w50_86),.acc(r50_86),.res(r50_87),.clk(clk),.wout(w50_87));
	PE pe50_88(.x(x88),.w(w50_87),.acc(r50_87),.res(r50_88),.clk(clk),.wout(w50_88));
	PE pe50_89(.x(x89),.w(w50_88),.acc(r50_88),.res(r50_89),.clk(clk),.wout(w50_89));
	PE pe50_90(.x(x90),.w(w50_89),.acc(r50_89),.res(r50_90),.clk(clk),.wout(w50_90));
	PE pe50_91(.x(x91),.w(w50_90),.acc(r50_90),.res(r50_91),.clk(clk),.wout(w50_91));
	PE pe50_92(.x(x92),.w(w50_91),.acc(r50_91),.res(r50_92),.clk(clk),.wout(w50_92));
	PE pe50_93(.x(x93),.w(w50_92),.acc(r50_92),.res(r50_93),.clk(clk),.wout(w50_93));
	PE pe50_94(.x(x94),.w(w50_93),.acc(r50_93),.res(r50_94),.clk(clk),.wout(w50_94));
	PE pe50_95(.x(x95),.w(w50_94),.acc(r50_94),.res(r50_95),.clk(clk),.wout(w50_95));
	PE pe50_96(.x(x96),.w(w50_95),.acc(r50_95),.res(r50_96),.clk(clk),.wout(w50_96));
	PE pe50_97(.x(x97),.w(w50_96),.acc(r50_96),.res(r50_97),.clk(clk),.wout(w50_97));
	PE pe50_98(.x(x98),.w(w50_97),.acc(r50_97),.res(r50_98),.clk(clk),.wout(w50_98));
	PE pe50_99(.x(x99),.w(w50_98),.acc(r50_98),.res(r50_99),.clk(clk),.wout(w50_99));
	PE pe50_100(.x(x100),.w(w50_99),.acc(r50_99),.res(r50_100),.clk(clk),.wout(w50_100));
	PE pe50_101(.x(x101),.w(w50_100),.acc(r50_100),.res(r50_101),.clk(clk),.wout(w50_101));
	PE pe50_102(.x(x102),.w(w50_101),.acc(r50_101),.res(r50_102),.clk(clk),.wout(w50_102));
	PE pe50_103(.x(x103),.w(w50_102),.acc(r50_102),.res(r50_103),.clk(clk),.wout(w50_103));
	PE pe50_104(.x(x104),.w(w50_103),.acc(r50_103),.res(r50_104),.clk(clk),.wout(w50_104));
	PE pe50_105(.x(x105),.w(w50_104),.acc(r50_104),.res(r50_105),.clk(clk),.wout(w50_105));
	PE pe50_106(.x(x106),.w(w50_105),.acc(r50_105),.res(r50_106),.clk(clk),.wout(w50_106));
	PE pe50_107(.x(x107),.w(w50_106),.acc(r50_106),.res(r50_107),.clk(clk),.wout(w50_107));
	PE pe50_108(.x(x108),.w(w50_107),.acc(r50_107),.res(r50_108),.clk(clk),.wout(w50_108));
	PE pe50_109(.x(x109),.w(w50_108),.acc(r50_108),.res(r50_109),.clk(clk),.wout(w50_109));
	PE pe50_110(.x(x110),.w(w50_109),.acc(r50_109),.res(r50_110),.clk(clk),.wout(w50_110));
	PE pe50_111(.x(x111),.w(w50_110),.acc(r50_110),.res(r50_111),.clk(clk),.wout(w50_111));
	PE pe50_112(.x(x112),.w(w50_111),.acc(r50_111),.res(r50_112),.clk(clk),.wout(w50_112));
	PE pe50_113(.x(x113),.w(w50_112),.acc(r50_112),.res(r50_113),.clk(clk),.wout(w50_113));
	PE pe50_114(.x(x114),.w(w50_113),.acc(r50_113),.res(r50_114),.clk(clk),.wout(w50_114));
	PE pe50_115(.x(x115),.w(w50_114),.acc(r50_114),.res(r50_115),.clk(clk),.wout(w50_115));
	PE pe50_116(.x(x116),.w(w50_115),.acc(r50_115),.res(r50_116),.clk(clk),.wout(w50_116));
	PE pe50_117(.x(x117),.w(w50_116),.acc(r50_116),.res(r50_117),.clk(clk),.wout(w50_117));
	PE pe50_118(.x(x118),.w(w50_117),.acc(r50_117),.res(r50_118),.clk(clk),.wout(w50_118));
	PE pe50_119(.x(x119),.w(w50_118),.acc(r50_118),.res(r50_119),.clk(clk),.wout(w50_119));
	PE pe50_120(.x(x120),.w(w50_119),.acc(r50_119),.res(r50_120),.clk(clk),.wout(w50_120));
	PE pe50_121(.x(x121),.w(w50_120),.acc(r50_120),.res(r50_121),.clk(clk),.wout(w50_121));
	PE pe50_122(.x(x122),.w(w50_121),.acc(r50_121),.res(r50_122),.clk(clk),.wout(w50_122));
	PE pe50_123(.x(x123),.w(w50_122),.acc(r50_122),.res(r50_123),.clk(clk),.wout(w50_123));
	PE pe50_124(.x(x124),.w(w50_123),.acc(r50_123),.res(r50_124),.clk(clk),.wout(w50_124));
	PE pe50_125(.x(x125),.w(w50_124),.acc(r50_124),.res(r50_125),.clk(clk),.wout(w50_125));
	PE pe50_126(.x(x126),.w(w50_125),.acc(r50_125),.res(r50_126),.clk(clk),.wout(w50_126));
	PE pe50_127(.x(x127),.w(w50_126),.acc(r50_126),.res(result50),.clk(clk),.wout(weight50));

	PE pe51_0(.x(x0),.w(w51),.acc(32'h0),.res(r51_0),.clk(clk),.wout(w51_0));
	PE pe51_1(.x(x1),.w(w51_0),.acc(r51_0),.res(r51_1),.clk(clk),.wout(w51_1));
	PE pe51_2(.x(x2),.w(w51_1),.acc(r51_1),.res(r51_2),.clk(clk),.wout(w51_2));
	PE pe51_3(.x(x3),.w(w51_2),.acc(r51_2),.res(r51_3),.clk(clk),.wout(w51_3));
	PE pe51_4(.x(x4),.w(w51_3),.acc(r51_3),.res(r51_4),.clk(clk),.wout(w51_4));
	PE pe51_5(.x(x5),.w(w51_4),.acc(r51_4),.res(r51_5),.clk(clk),.wout(w51_5));
	PE pe51_6(.x(x6),.w(w51_5),.acc(r51_5),.res(r51_6),.clk(clk),.wout(w51_6));
	PE pe51_7(.x(x7),.w(w51_6),.acc(r51_6),.res(r51_7),.clk(clk),.wout(w51_7));
	PE pe51_8(.x(x8),.w(w51_7),.acc(r51_7),.res(r51_8),.clk(clk),.wout(w51_8));
	PE pe51_9(.x(x9),.w(w51_8),.acc(r51_8),.res(r51_9),.clk(clk),.wout(w51_9));
	PE pe51_10(.x(x10),.w(w51_9),.acc(r51_9),.res(r51_10),.clk(clk),.wout(w51_10));
	PE pe51_11(.x(x11),.w(w51_10),.acc(r51_10),.res(r51_11),.clk(clk),.wout(w51_11));
	PE pe51_12(.x(x12),.w(w51_11),.acc(r51_11),.res(r51_12),.clk(clk),.wout(w51_12));
	PE pe51_13(.x(x13),.w(w51_12),.acc(r51_12),.res(r51_13),.clk(clk),.wout(w51_13));
	PE pe51_14(.x(x14),.w(w51_13),.acc(r51_13),.res(r51_14),.clk(clk),.wout(w51_14));
	PE pe51_15(.x(x15),.w(w51_14),.acc(r51_14),.res(r51_15),.clk(clk),.wout(w51_15));
	PE pe51_16(.x(x16),.w(w51_15),.acc(r51_15),.res(r51_16),.clk(clk),.wout(w51_16));
	PE pe51_17(.x(x17),.w(w51_16),.acc(r51_16),.res(r51_17),.clk(clk),.wout(w51_17));
	PE pe51_18(.x(x18),.w(w51_17),.acc(r51_17),.res(r51_18),.clk(clk),.wout(w51_18));
	PE pe51_19(.x(x19),.w(w51_18),.acc(r51_18),.res(r51_19),.clk(clk),.wout(w51_19));
	PE pe51_20(.x(x20),.w(w51_19),.acc(r51_19),.res(r51_20),.clk(clk),.wout(w51_20));
	PE pe51_21(.x(x21),.w(w51_20),.acc(r51_20),.res(r51_21),.clk(clk),.wout(w51_21));
	PE pe51_22(.x(x22),.w(w51_21),.acc(r51_21),.res(r51_22),.clk(clk),.wout(w51_22));
	PE pe51_23(.x(x23),.w(w51_22),.acc(r51_22),.res(r51_23),.clk(clk),.wout(w51_23));
	PE pe51_24(.x(x24),.w(w51_23),.acc(r51_23),.res(r51_24),.clk(clk),.wout(w51_24));
	PE pe51_25(.x(x25),.w(w51_24),.acc(r51_24),.res(r51_25),.clk(clk),.wout(w51_25));
	PE pe51_26(.x(x26),.w(w51_25),.acc(r51_25),.res(r51_26),.clk(clk),.wout(w51_26));
	PE pe51_27(.x(x27),.w(w51_26),.acc(r51_26),.res(r51_27),.clk(clk),.wout(w51_27));
	PE pe51_28(.x(x28),.w(w51_27),.acc(r51_27),.res(r51_28),.clk(clk),.wout(w51_28));
	PE pe51_29(.x(x29),.w(w51_28),.acc(r51_28),.res(r51_29),.clk(clk),.wout(w51_29));
	PE pe51_30(.x(x30),.w(w51_29),.acc(r51_29),.res(r51_30),.clk(clk),.wout(w51_30));
	PE pe51_31(.x(x31),.w(w51_30),.acc(r51_30),.res(r51_31),.clk(clk),.wout(w51_31));
	PE pe51_32(.x(x32),.w(w51_31),.acc(r51_31),.res(r51_32),.clk(clk),.wout(w51_32));
	PE pe51_33(.x(x33),.w(w51_32),.acc(r51_32),.res(r51_33),.clk(clk),.wout(w51_33));
	PE pe51_34(.x(x34),.w(w51_33),.acc(r51_33),.res(r51_34),.clk(clk),.wout(w51_34));
	PE pe51_35(.x(x35),.w(w51_34),.acc(r51_34),.res(r51_35),.clk(clk),.wout(w51_35));
	PE pe51_36(.x(x36),.w(w51_35),.acc(r51_35),.res(r51_36),.clk(clk),.wout(w51_36));
	PE pe51_37(.x(x37),.w(w51_36),.acc(r51_36),.res(r51_37),.clk(clk),.wout(w51_37));
	PE pe51_38(.x(x38),.w(w51_37),.acc(r51_37),.res(r51_38),.clk(clk),.wout(w51_38));
	PE pe51_39(.x(x39),.w(w51_38),.acc(r51_38),.res(r51_39),.clk(clk),.wout(w51_39));
	PE pe51_40(.x(x40),.w(w51_39),.acc(r51_39),.res(r51_40),.clk(clk),.wout(w51_40));
	PE pe51_41(.x(x41),.w(w51_40),.acc(r51_40),.res(r51_41),.clk(clk),.wout(w51_41));
	PE pe51_42(.x(x42),.w(w51_41),.acc(r51_41),.res(r51_42),.clk(clk),.wout(w51_42));
	PE pe51_43(.x(x43),.w(w51_42),.acc(r51_42),.res(r51_43),.clk(clk),.wout(w51_43));
	PE pe51_44(.x(x44),.w(w51_43),.acc(r51_43),.res(r51_44),.clk(clk),.wout(w51_44));
	PE pe51_45(.x(x45),.w(w51_44),.acc(r51_44),.res(r51_45),.clk(clk),.wout(w51_45));
	PE pe51_46(.x(x46),.w(w51_45),.acc(r51_45),.res(r51_46),.clk(clk),.wout(w51_46));
	PE pe51_47(.x(x47),.w(w51_46),.acc(r51_46),.res(r51_47),.clk(clk),.wout(w51_47));
	PE pe51_48(.x(x48),.w(w51_47),.acc(r51_47),.res(r51_48),.clk(clk),.wout(w51_48));
	PE pe51_49(.x(x49),.w(w51_48),.acc(r51_48),.res(r51_49),.clk(clk),.wout(w51_49));
	PE pe51_50(.x(x50),.w(w51_49),.acc(r51_49),.res(r51_50),.clk(clk),.wout(w51_50));
	PE pe51_51(.x(x51),.w(w51_50),.acc(r51_50),.res(r51_51),.clk(clk),.wout(w51_51));
	PE pe51_52(.x(x52),.w(w51_51),.acc(r51_51),.res(r51_52),.clk(clk),.wout(w51_52));
	PE pe51_53(.x(x53),.w(w51_52),.acc(r51_52),.res(r51_53),.clk(clk),.wout(w51_53));
	PE pe51_54(.x(x54),.w(w51_53),.acc(r51_53),.res(r51_54),.clk(clk),.wout(w51_54));
	PE pe51_55(.x(x55),.w(w51_54),.acc(r51_54),.res(r51_55),.clk(clk),.wout(w51_55));
	PE pe51_56(.x(x56),.w(w51_55),.acc(r51_55),.res(r51_56),.clk(clk),.wout(w51_56));
	PE pe51_57(.x(x57),.w(w51_56),.acc(r51_56),.res(r51_57),.clk(clk),.wout(w51_57));
	PE pe51_58(.x(x58),.w(w51_57),.acc(r51_57),.res(r51_58),.clk(clk),.wout(w51_58));
	PE pe51_59(.x(x59),.w(w51_58),.acc(r51_58),.res(r51_59),.clk(clk),.wout(w51_59));
	PE pe51_60(.x(x60),.w(w51_59),.acc(r51_59),.res(r51_60),.clk(clk),.wout(w51_60));
	PE pe51_61(.x(x61),.w(w51_60),.acc(r51_60),.res(r51_61),.clk(clk),.wout(w51_61));
	PE pe51_62(.x(x62),.w(w51_61),.acc(r51_61),.res(r51_62),.clk(clk),.wout(w51_62));
	PE pe51_63(.x(x63),.w(w51_62),.acc(r51_62),.res(r51_63),.clk(clk),.wout(w51_63));
	PE pe51_64(.x(x64),.w(w51_63),.acc(r51_63),.res(r51_64),.clk(clk),.wout(w51_64));
	PE pe51_65(.x(x65),.w(w51_64),.acc(r51_64),.res(r51_65),.clk(clk),.wout(w51_65));
	PE pe51_66(.x(x66),.w(w51_65),.acc(r51_65),.res(r51_66),.clk(clk),.wout(w51_66));
	PE pe51_67(.x(x67),.w(w51_66),.acc(r51_66),.res(r51_67),.clk(clk),.wout(w51_67));
	PE pe51_68(.x(x68),.w(w51_67),.acc(r51_67),.res(r51_68),.clk(clk),.wout(w51_68));
	PE pe51_69(.x(x69),.w(w51_68),.acc(r51_68),.res(r51_69),.clk(clk),.wout(w51_69));
	PE pe51_70(.x(x70),.w(w51_69),.acc(r51_69),.res(r51_70),.clk(clk),.wout(w51_70));
	PE pe51_71(.x(x71),.w(w51_70),.acc(r51_70),.res(r51_71),.clk(clk),.wout(w51_71));
	PE pe51_72(.x(x72),.w(w51_71),.acc(r51_71),.res(r51_72),.clk(clk),.wout(w51_72));
	PE pe51_73(.x(x73),.w(w51_72),.acc(r51_72),.res(r51_73),.clk(clk),.wout(w51_73));
	PE pe51_74(.x(x74),.w(w51_73),.acc(r51_73),.res(r51_74),.clk(clk),.wout(w51_74));
	PE pe51_75(.x(x75),.w(w51_74),.acc(r51_74),.res(r51_75),.clk(clk),.wout(w51_75));
	PE pe51_76(.x(x76),.w(w51_75),.acc(r51_75),.res(r51_76),.clk(clk),.wout(w51_76));
	PE pe51_77(.x(x77),.w(w51_76),.acc(r51_76),.res(r51_77),.clk(clk),.wout(w51_77));
	PE pe51_78(.x(x78),.w(w51_77),.acc(r51_77),.res(r51_78),.clk(clk),.wout(w51_78));
	PE pe51_79(.x(x79),.w(w51_78),.acc(r51_78),.res(r51_79),.clk(clk),.wout(w51_79));
	PE pe51_80(.x(x80),.w(w51_79),.acc(r51_79),.res(r51_80),.clk(clk),.wout(w51_80));
	PE pe51_81(.x(x81),.w(w51_80),.acc(r51_80),.res(r51_81),.clk(clk),.wout(w51_81));
	PE pe51_82(.x(x82),.w(w51_81),.acc(r51_81),.res(r51_82),.clk(clk),.wout(w51_82));
	PE pe51_83(.x(x83),.w(w51_82),.acc(r51_82),.res(r51_83),.clk(clk),.wout(w51_83));
	PE pe51_84(.x(x84),.w(w51_83),.acc(r51_83),.res(r51_84),.clk(clk),.wout(w51_84));
	PE pe51_85(.x(x85),.w(w51_84),.acc(r51_84),.res(r51_85),.clk(clk),.wout(w51_85));
	PE pe51_86(.x(x86),.w(w51_85),.acc(r51_85),.res(r51_86),.clk(clk),.wout(w51_86));
	PE pe51_87(.x(x87),.w(w51_86),.acc(r51_86),.res(r51_87),.clk(clk),.wout(w51_87));
	PE pe51_88(.x(x88),.w(w51_87),.acc(r51_87),.res(r51_88),.clk(clk),.wout(w51_88));
	PE pe51_89(.x(x89),.w(w51_88),.acc(r51_88),.res(r51_89),.clk(clk),.wout(w51_89));
	PE pe51_90(.x(x90),.w(w51_89),.acc(r51_89),.res(r51_90),.clk(clk),.wout(w51_90));
	PE pe51_91(.x(x91),.w(w51_90),.acc(r51_90),.res(r51_91),.clk(clk),.wout(w51_91));
	PE pe51_92(.x(x92),.w(w51_91),.acc(r51_91),.res(r51_92),.clk(clk),.wout(w51_92));
	PE pe51_93(.x(x93),.w(w51_92),.acc(r51_92),.res(r51_93),.clk(clk),.wout(w51_93));
	PE pe51_94(.x(x94),.w(w51_93),.acc(r51_93),.res(r51_94),.clk(clk),.wout(w51_94));
	PE pe51_95(.x(x95),.w(w51_94),.acc(r51_94),.res(r51_95),.clk(clk),.wout(w51_95));
	PE pe51_96(.x(x96),.w(w51_95),.acc(r51_95),.res(r51_96),.clk(clk),.wout(w51_96));
	PE pe51_97(.x(x97),.w(w51_96),.acc(r51_96),.res(r51_97),.clk(clk),.wout(w51_97));
	PE pe51_98(.x(x98),.w(w51_97),.acc(r51_97),.res(r51_98),.clk(clk),.wout(w51_98));
	PE pe51_99(.x(x99),.w(w51_98),.acc(r51_98),.res(r51_99),.clk(clk),.wout(w51_99));
	PE pe51_100(.x(x100),.w(w51_99),.acc(r51_99),.res(r51_100),.clk(clk),.wout(w51_100));
	PE pe51_101(.x(x101),.w(w51_100),.acc(r51_100),.res(r51_101),.clk(clk),.wout(w51_101));
	PE pe51_102(.x(x102),.w(w51_101),.acc(r51_101),.res(r51_102),.clk(clk),.wout(w51_102));
	PE pe51_103(.x(x103),.w(w51_102),.acc(r51_102),.res(r51_103),.clk(clk),.wout(w51_103));
	PE pe51_104(.x(x104),.w(w51_103),.acc(r51_103),.res(r51_104),.clk(clk),.wout(w51_104));
	PE pe51_105(.x(x105),.w(w51_104),.acc(r51_104),.res(r51_105),.clk(clk),.wout(w51_105));
	PE pe51_106(.x(x106),.w(w51_105),.acc(r51_105),.res(r51_106),.clk(clk),.wout(w51_106));
	PE pe51_107(.x(x107),.w(w51_106),.acc(r51_106),.res(r51_107),.clk(clk),.wout(w51_107));
	PE pe51_108(.x(x108),.w(w51_107),.acc(r51_107),.res(r51_108),.clk(clk),.wout(w51_108));
	PE pe51_109(.x(x109),.w(w51_108),.acc(r51_108),.res(r51_109),.clk(clk),.wout(w51_109));
	PE pe51_110(.x(x110),.w(w51_109),.acc(r51_109),.res(r51_110),.clk(clk),.wout(w51_110));
	PE pe51_111(.x(x111),.w(w51_110),.acc(r51_110),.res(r51_111),.clk(clk),.wout(w51_111));
	PE pe51_112(.x(x112),.w(w51_111),.acc(r51_111),.res(r51_112),.clk(clk),.wout(w51_112));
	PE pe51_113(.x(x113),.w(w51_112),.acc(r51_112),.res(r51_113),.clk(clk),.wout(w51_113));
	PE pe51_114(.x(x114),.w(w51_113),.acc(r51_113),.res(r51_114),.clk(clk),.wout(w51_114));
	PE pe51_115(.x(x115),.w(w51_114),.acc(r51_114),.res(r51_115),.clk(clk),.wout(w51_115));
	PE pe51_116(.x(x116),.w(w51_115),.acc(r51_115),.res(r51_116),.clk(clk),.wout(w51_116));
	PE pe51_117(.x(x117),.w(w51_116),.acc(r51_116),.res(r51_117),.clk(clk),.wout(w51_117));
	PE pe51_118(.x(x118),.w(w51_117),.acc(r51_117),.res(r51_118),.clk(clk),.wout(w51_118));
	PE pe51_119(.x(x119),.w(w51_118),.acc(r51_118),.res(r51_119),.clk(clk),.wout(w51_119));
	PE pe51_120(.x(x120),.w(w51_119),.acc(r51_119),.res(r51_120),.clk(clk),.wout(w51_120));
	PE pe51_121(.x(x121),.w(w51_120),.acc(r51_120),.res(r51_121),.clk(clk),.wout(w51_121));
	PE pe51_122(.x(x122),.w(w51_121),.acc(r51_121),.res(r51_122),.clk(clk),.wout(w51_122));
	PE pe51_123(.x(x123),.w(w51_122),.acc(r51_122),.res(r51_123),.clk(clk),.wout(w51_123));
	PE pe51_124(.x(x124),.w(w51_123),.acc(r51_123),.res(r51_124),.clk(clk),.wout(w51_124));
	PE pe51_125(.x(x125),.w(w51_124),.acc(r51_124),.res(r51_125),.clk(clk),.wout(w51_125));
	PE pe51_126(.x(x126),.w(w51_125),.acc(r51_125),.res(r51_126),.clk(clk),.wout(w51_126));
	PE pe51_127(.x(x127),.w(w51_126),.acc(r51_126),.res(result51),.clk(clk),.wout(weight51));

	PE pe52_0(.x(x0),.w(w52),.acc(32'h0),.res(r52_0),.clk(clk),.wout(w52_0));
	PE pe52_1(.x(x1),.w(w52_0),.acc(r52_0),.res(r52_1),.clk(clk),.wout(w52_1));
	PE pe52_2(.x(x2),.w(w52_1),.acc(r52_1),.res(r52_2),.clk(clk),.wout(w52_2));
	PE pe52_3(.x(x3),.w(w52_2),.acc(r52_2),.res(r52_3),.clk(clk),.wout(w52_3));
	PE pe52_4(.x(x4),.w(w52_3),.acc(r52_3),.res(r52_4),.clk(clk),.wout(w52_4));
	PE pe52_5(.x(x5),.w(w52_4),.acc(r52_4),.res(r52_5),.clk(clk),.wout(w52_5));
	PE pe52_6(.x(x6),.w(w52_5),.acc(r52_5),.res(r52_6),.clk(clk),.wout(w52_6));
	PE pe52_7(.x(x7),.w(w52_6),.acc(r52_6),.res(r52_7),.clk(clk),.wout(w52_7));
	PE pe52_8(.x(x8),.w(w52_7),.acc(r52_7),.res(r52_8),.clk(clk),.wout(w52_8));
	PE pe52_9(.x(x9),.w(w52_8),.acc(r52_8),.res(r52_9),.clk(clk),.wout(w52_9));
	PE pe52_10(.x(x10),.w(w52_9),.acc(r52_9),.res(r52_10),.clk(clk),.wout(w52_10));
	PE pe52_11(.x(x11),.w(w52_10),.acc(r52_10),.res(r52_11),.clk(clk),.wout(w52_11));
	PE pe52_12(.x(x12),.w(w52_11),.acc(r52_11),.res(r52_12),.clk(clk),.wout(w52_12));
	PE pe52_13(.x(x13),.w(w52_12),.acc(r52_12),.res(r52_13),.clk(clk),.wout(w52_13));
	PE pe52_14(.x(x14),.w(w52_13),.acc(r52_13),.res(r52_14),.clk(clk),.wout(w52_14));
	PE pe52_15(.x(x15),.w(w52_14),.acc(r52_14),.res(r52_15),.clk(clk),.wout(w52_15));
	PE pe52_16(.x(x16),.w(w52_15),.acc(r52_15),.res(r52_16),.clk(clk),.wout(w52_16));
	PE pe52_17(.x(x17),.w(w52_16),.acc(r52_16),.res(r52_17),.clk(clk),.wout(w52_17));
	PE pe52_18(.x(x18),.w(w52_17),.acc(r52_17),.res(r52_18),.clk(clk),.wout(w52_18));
	PE pe52_19(.x(x19),.w(w52_18),.acc(r52_18),.res(r52_19),.clk(clk),.wout(w52_19));
	PE pe52_20(.x(x20),.w(w52_19),.acc(r52_19),.res(r52_20),.clk(clk),.wout(w52_20));
	PE pe52_21(.x(x21),.w(w52_20),.acc(r52_20),.res(r52_21),.clk(clk),.wout(w52_21));
	PE pe52_22(.x(x22),.w(w52_21),.acc(r52_21),.res(r52_22),.clk(clk),.wout(w52_22));
	PE pe52_23(.x(x23),.w(w52_22),.acc(r52_22),.res(r52_23),.clk(clk),.wout(w52_23));
	PE pe52_24(.x(x24),.w(w52_23),.acc(r52_23),.res(r52_24),.clk(clk),.wout(w52_24));
	PE pe52_25(.x(x25),.w(w52_24),.acc(r52_24),.res(r52_25),.clk(clk),.wout(w52_25));
	PE pe52_26(.x(x26),.w(w52_25),.acc(r52_25),.res(r52_26),.clk(clk),.wout(w52_26));
	PE pe52_27(.x(x27),.w(w52_26),.acc(r52_26),.res(r52_27),.clk(clk),.wout(w52_27));
	PE pe52_28(.x(x28),.w(w52_27),.acc(r52_27),.res(r52_28),.clk(clk),.wout(w52_28));
	PE pe52_29(.x(x29),.w(w52_28),.acc(r52_28),.res(r52_29),.clk(clk),.wout(w52_29));
	PE pe52_30(.x(x30),.w(w52_29),.acc(r52_29),.res(r52_30),.clk(clk),.wout(w52_30));
	PE pe52_31(.x(x31),.w(w52_30),.acc(r52_30),.res(r52_31),.clk(clk),.wout(w52_31));
	PE pe52_32(.x(x32),.w(w52_31),.acc(r52_31),.res(r52_32),.clk(clk),.wout(w52_32));
	PE pe52_33(.x(x33),.w(w52_32),.acc(r52_32),.res(r52_33),.clk(clk),.wout(w52_33));
	PE pe52_34(.x(x34),.w(w52_33),.acc(r52_33),.res(r52_34),.clk(clk),.wout(w52_34));
	PE pe52_35(.x(x35),.w(w52_34),.acc(r52_34),.res(r52_35),.clk(clk),.wout(w52_35));
	PE pe52_36(.x(x36),.w(w52_35),.acc(r52_35),.res(r52_36),.clk(clk),.wout(w52_36));
	PE pe52_37(.x(x37),.w(w52_36),.acc(r52_36),.res(r52_37),.clk(clk),.wout(w52_37));
	PE pe52_38(.x(x38),.w(w52_37),.acc(r52_37),.res(r52_38),.clk(clk),.wout(w52_38));
	PE pe52_39(.x(x39),.w(w52_38),.acc(r52_38),.res(r52_39),.clk(clk),.wout(w52_39));
	PE pe52_40(.x(x40),.w(w52_39),.acc(r52_39),.res(r52_40),.clk(clk),.wout(w52_40));
	PE pe52_41(.x(x41),.w(w52_40),.acc(r52_40),.res(r52_41),.clk(clk),.wout(w52_41));
	PE pe52_42(.x(x42),.w(w52_41),.acc(r52_41),.res(r52_42),.clk(clk),.wout(w52_42));
	PE pe52_43(.x(x43),.w(w52_42),.acc(r52_42),.res(r52_43),.clk(clk),.wout(w52_43));
	PE pe52_44(.x(x44),.w(w52_43),.acc(r52_43),.res(r52_44),.clk(clk),.wout(w52_44));
	PE pe52_45(.x(x45),.w(w52_44),.acc(r52_44),.res(r52_45),.clk(clk),.wout(w52_45));
	PE pe52_46(.x(x46),.w(w52_45),.acc(r52_45),.res(r52_46),.clk(clk),.wout(w52_46));
	PE pe52_47(.x(x47),.w(w52_46),.acc(r52_46),.res(r52_47),.clk(clk),.wout(w52_47));
	PE pe52_48(.x(x48),.w(w52_47),.acc(r52_47),.res(r52_48),.clk(clk),.wout(w52_48));
	PE pe52_49(.x(x49),.w(w52_48),.acc(r52_48),.res(r52_49),.clk(clk),.wout(w52_49));
	PE pe52_50(.x(x50),.w(w52_49),.acc(r52_49),.res(r52_50),.clk(clk),.wout(w52_50));
	PE pe52_51(.x(x51),.w(w52_50),.acc(r52_50),.res(r52_51),.clk(clk),.wout(w52_51));
	PE pe52_52(.x(x52),.w(w52_51),.acc(r52_51),.res(r52_52),.clk(clk),.wout(w52_52));
	PE pe52_53(.x(x53),.w(w52_52),.acc(r52_52),.res(r52_53),.clk(clk),.wout(w52_53));
	PE pe52_54(.x(x54),.w(w52_53),.acc(r52_53),.res(r52_54),.clk(clk),.wout(w52_54));
	PE pe52_55(.x(x55),.w(w52_54),.acc(r52_54),.res(r52_55),.clk(clk),.wout(w52_55));
	PE pe52_56(.x(x56),.w(w52_55),.acc(r52_55),.res(r52_56),.clk(clk),.wout(w52_56));
	PE pe52_57(.x(x57),.w(w52_56),.acc(r52_56),.res(r52_57),.clk(clk),.wout(w52_57));
	PE pe52_58(.x(x58),.w(w52_57),.acc(r52_57),.res(r52_58),.clk(clk),.wout(w52_58));
	PE pe52_59(.x(x59),.w(w52_58),.acc(r52_58),.res(r52_59),.clk(clk),.wout(w52_59));
	PE pe52_60(.x(x60),.w(w52_59),.acc(r52_59),.res(r52_60),.clk(clk),.wout(w52_60));
	PE pe52_61(.x(x61),.w(w52_60),.acc(r52_60),.res(r52_61),.clk(clk),.wout(w52_61));
	PE pe52_62(.x(x62),.w(w52_61),.acc(r52_61),.res(r52_62),.clk(clk),.wout(w52_62));
	PE pe52_63(.x(x63),.w(w52_62),.acc(r52_62),.res(r52_63),.clk(clk),.wout(w52_63));
	PE pe52_64(.x(x64),.w(w52_63),.acc(r52_63),.res(r52_64),.clk(clk),.wout(w52_64));
	PE pe52_65(.x(x65),.w(w52_64),.acc(r52_64),.res(r52_65),.clk(clk),.wout(w52_65));
	PE pe52_66(.x(x66),.w(w52_65),.acc(r52_65),.res(r52_66),.clk(clk),.wout(w52_66));
	PE pe52_67(.x(x67),.w(w52_66),.acc(r52_66),.res(r52_67),.clk(clk),.wout(w52_67));
	PE pe52_68(.x(x68),.w(w52_67),.acc(r52_67),.res(r52_68),.clk(clk),.wout(w52_68));
	PE pe52_69(.x(x69),.w(w52_68),.acc(r52_68),.res(r52_69),.clk(clk),.wout(w52_69));
	PE pe52_70(.x(x70),.w(w52_69),.acc(r52_69),.res(r52_70),.clk(clk),.wout(w52_70));
	PE pe52_71(.x(x71),.w(w52_70),.acc(r52_70),.res(r52_71),.clk(clk),.wout(w52_71));
	PE pe52_72(.x(x72),.w(w52_71),.acc(r52_71),.res(r52_72),.clk(clk),.wout(w52_72));
	PE pe52_73(.x(x73),.w(w52_72),.acc(r52_72),.res(r52_73),.clk(clk),.wout(w52_73));
	PE pe52_74(.x(x74),.w(w52_73),.acc(r52_73),.res(r52_74),.clk(clk),.wout(w52_74));
	PE pe52_75(.x(x75),.w(w52_74),.acc(r52_74),.res(r52_75),.clk(clk),.wout(w52_75));
	PE pe52_76(.x(x76),.w(w52_75),.acc(r52_75),.res(r52_76),.clk(clk),.wout(w52_76));
	PE pe52_77(.x(x77),.w(w52_76),.acc(r52_76),.res(r52_77),.clk(clk),.wout(w52_77));
	PE pe52_78(.x(x78),.w(w52_77),.acc(r52_77),.res(r52_78),.clk(clk),.wout(w52_78));
	PE pe52_79(.x(x79),.w(w52_78),.acc(r52_78),.res(r52_79),.clk(clk),.wout(w52_79));
	PE pe52_80(.x(x80),.w(w52_79),.acc(r52_79),.res(r52_80),.clk(clk),.wout(w52_80));
	PE pe52_81(.x(x81),.w(w52_80),.acc(r52_80),.res(r52_81),.clk(clk),.wout(w52_81));
	PE pe52_82(.x(x82),.w(w52_81),.acc(r52_81),.res(r52_82),.clk(clk),.wout(w52_82));
	PE pe52_83(.x(x83),.w(w52_82),.acc(r52_82),.res(r52_83),.clk(clk),.wout(w52_83));
	PE pe52_84(.x(x84),.w(w52_83),.acc(r52_83),.res(r52_84),.clk(clk),.wout(w52_84));
	PE pe52_85(.x(x85),.w(w52_84),.acc(r52_84),.res(r52_85),.clk(clk),.wout(w52_85));
	PE pe52_86(.x(x86),.w(w52_85),.acc(r52_85),.res(r52_86),.clk(clk),.wout(w52_86));
	PE pe52_87(.x(x87),.w(w52_86),.acc(r52_86),.res(r52_87),.clk(clk),.wout(w52_87));
	PE pe52_88(.x(x88),.w(w52_87),.acc(r52_87),.res(r52_88),.clk(clk),.wout(w52_88));
	PE pe52_89(.x(x89),.w(w52_88),.acc(r52_88),.res(r52_89),.clk(clk),.wout(w52_89));
	PE pe52_90(.x(x90),.w(w52_89),.acc(r52_89),.res(r52_90),.clk(clk),.wout(w52_90));
	PE pe52_91(.x(x91),.w(w52_90),.acc(r52_90),.res(r52_91),.clk(clk),.wout(w52_91));
	PE pe52_92(.x(x92),.w(w52_91),.acc(r52_91),.res(r52_92),.clk(clk),.wout(w52_92));
	PE pe52_93(.x(x93),.w(w52_92),.acc(r52_92),.res(r52_93),.clk(clk),.wout(w52_93));
	PE pe52_94(.x(x94),.w(w52_93),.acc(r52_93),.res(r52_94),.clk(clk),.wout(w52_94));
	PE pe52_95(.x(x95),.w(w52_94),.acc(r52_94),.res(r52_95),.clk(clk),.wout(w52_95));
	PE pe52_96(.x(x96),.w(w52_95),.acc(r52_95),.res(r52_96),.clk(clk),.wout(w52_96));
	PE pe52_97(.x(x97),.w(w52_96),.acc(r52_96),.res(r52_97),.clk(clk),.wout(w52_97));
	PE pe52_98(.x(x98),.w(w52_97),.acc(r52_97),.res(r52_98),.clk(clk),.wout(w52_98));
	PE pe52_99(.x(x99),.w(w52_98),.acc(r52_98),.res(r52_99),.clk(clk),.wout(w52_99));
	PE pe52_100(.x(x100),.w(w52_99),.acc(r52_99),.res(r52_100),.clk(clk),.wout(w52_100));
	PE pe52_101(.x(x101),.w(w52_100),.acc(r52_100),.res(r52_101),.clk(clk),.wout(w52_101));
	PE pe52_102(.x(x102),.w(w52_101),.acc(r52_101),.res(r52_102),.clk(clk),.wout(w52_102));
	PE pe52_103(.x(x103),.w(w52_102),.acc(r52_102),.res(r52_103),.clk(clk),.wout(w52_103));
	PE pe52_104(.x(x104),.w(w52_103),.acc(r52_103),.res(r52_104),.clk(clk),.wout(w52_104));
	PE pe52_105(.x(x105),.w(w52_104),.acc(r52_104),.res(r52_105),.clk(clk),.wout(w52_105));
	PE pe52_106(.x(x106),.w(w52_105),.acc(r52_105),.res(r52_106),.clk(clk),.wout(w52_106));
	PE pe52_107(.x(x107),.w(w52_106),.acc(r52_106),.res(r52_107),.clk(clk),.wout(w52_107));
	PE pe52_108(.x(x108),.w(w52_107),.acc(r52_107),.res(r52_108),.clk(clk),.wout(w52_108));
	PE pe52_109(.x(x109),.w(w52_108),.acc(r52_108),.res(r52_109),.clk(clk),.wout(w52_109));
	PE pe52_110(.x(x110),.w(w52_109),.acc(r52_109),.res(r52_110),.clk(clk),.wout(w52_110));
	PE pe52_111(.x(x111),.w(w52_110),.acc(r52_110),.res(r52_111),.clk(clk),.wout(w52_111));
	PE pe52_112(.x(x112),.w(w52_111),.acc(r52_111),.res(r52_112),.clk(clk),.wout(w52_112));
	PE pe52_113(.x(x113),.w(w52_112),.acc(r52_112),.res(r52_113),.clk(clk),.wout(w52_113));
	PE pe52_114(.x(x114),.w(w52_113),.acc(r52_113),.res(r52_114),.clk(clk),.wout(w52_114));
	PE pe52_115(.x(x115),.w(w52_114),.acc(r52_114),.res(r52_115),.clk(clk),.wout(w52_115));
	PE pe52_116(.x(x116),.w(w52_115),.acc(r52_115),.res(r52_116),.clk(clk),.wout(w52_116));
	PE pe52_117(.x(x117),.w(w52_116),.acc(r52_116),.res(r52_117),.clk(clk),.wout(w52_117));
	PE pe52_118(.x(x118),.w(w52_117),.acc(r52_117),.res(r52_118),.clk(clk),.wout(w52_118));
	PE pe52_119(.x(x119),.w(w52_118),.acc(r52_118),.res(r52_119),.clk(clk),.wout(w52_119));
	PE pe52_120(.x(x120),.w(w52_119),.acc(r52_119),.res(r52_120),.clk(clk),.wout(w52_120));
	PE pe52_121(.x(x121),.w(w52_120),.acc(r52_120),.res(r52_121),.clk(clk),.wout(w52_121));
	PE pe52_122(.x(x122),.w(w52_121),.acc(r52_121),.res(r52_122),.clk(clk),.wout(w52_122));
	PE pe52_123(.x(x123),.w(w52_122),.acc(r52_122),.res(r52_123),.clk(clk),.wout(w52_123));
	PE pe52_124(.x(x124),.w(w52_123),.acc(r52_123),.res(r52_124),.clk(clk),.wout(w52_124));
	PE pe52_125(.x(x125),.w(w52_124),.acc(r52_124),.res(r52_125),.clk(clk),.wout(w52_125));
	PE pe52_126(.x(x126),.w(w52_125),.acc(r52_125),.res(r52_126),.clk(clk),.wout(w52_126));
	PE pe52_127(.x(x127),.w(w52_126),.acc(r52_126),.res(result52),.clk(clk),.wout(weight52));

	PE pe53_0(.x(x0),.w(w53),.acc(32'h0),.res(r53_0),.clk(clk),.wout(w53_0));
	PE pe53_1(.x(x1),.w(w53_0),.acc(r53_0),.res(r53_1),.clk(clk),.wout(w53_1));
	PE pe53_2(.x(x2),.w(w53_1),.acc(r53_1),.res(r53_2),.clk(clk),.wout(w53_2));
	PE pe53_3(.x(x3),.w(w53_2),.acc(r53_2),.res(r53_3),.clk(clk),.wout(w53_3));
	PE pe53_4(.x(x4),.w(w53_3),.acc(r53_3),.res(r53_4),.clk(clk),.wout(w53_4));
	PE pe53_5(.x(x5),.w(w53_4),.acc(r53_4),.res(r53_5),.clk(clk),.wout(w53_5));
	PE pe53_6(.x(x6),.w(w53_5),.acc(r53_5),.res(r53_6),.clk(clk),.wout(w53_6));
	PE pe53_7(.x(x7),.w(w53_6),.acc(r53_6),.res(r53_7),.clk(clk),.wout(w53_7));
	PE pe53_8(.x(x8),.w(w53_7),.acc(r53_7),.res(r53_8),.clk(clk),.wout(w53_8));
	PE pe53_9(.x(x9),.w(w53_8),.acc(r53_8),.res(r53_9),.clk(clk),.wout(w53_9));
	PE pe53_10(.x(x10),.w(w53_9),.acc(r53_9),.res(r53_10),.clk(clk),.wout(w53_10));
	PE pe53_11(.x(x11),.w(w53_10),.acc(r53_10),.res(r53_11),.clk(clk),.wout(w53_11));
	PE pe53_12(.x(x12),.w(w53_11),.acc(r53_11),.res(r53_12),.clk(clk),.wout(w53_12));
	PE pe53_13(.x(x13),.w(w53_12),.acc(r53_12),.res(r53_13),.clk(clk),.wout(w53_13));
	PE pe53_14(.x(x14),.w(w53_13),.acc(r53_13),.res(r53_14),.clk(clk),.wout(w53_14));
	PE pe53_15(.x(x15),.w(w53_14),.acc(r53_14),.res(r53_15),.clk(clk),.wout(w53_15));
	PE pe53_16(.x(x16),.w(w53_15),.acc(r53_15),.res(r53_16),.clk(clk),.wout(w53_16));
	PE pe53_17(.x(x17),.w(w53_16),.acc(r53_16),.res(r53_17),.clk(clk),.wout(w53_17));
	PE pe53_18(.x(x18),.w(w53_17),.acc(r53_17),.res(r53_18),.clk(clk),.wout(w53_18));
	PE pe53_19(.x(x19),.w(w53_18),.acc(r53_18),.res(r53_19),.clk(clk),.wout(w53_19));
	PE pe53_20(.x(x20),.w(w53_19),.acc(r53_19),.res(r53_20),.clk(clk),.wout(w53_20));
	PE pe53_21(.x(x21),.w(w53_20),.acc(r53_20),.res(r53_21),.clk(clk),.wout(w53_21));
	PE pe53_22(.x(x22),.w(w53_21),.acc(r53_21),.res(r53_22),.clk(clk),.wout(w53_22));
	PE pe53_23(.x(x23),.w(w53_22),.acc(r53_22),.res(r53_23),.clk(clk),.wout(w53_23));
	PE pe53_24(.x(x24),.w(w53_23),.acc(r53_23),.res(r53_24),.clk(clk),.wout(w53_24));
	PE pe53_25(.x(x25),.w(w53_24),.acc(r53_24),.res(r53_25),.clk(clk),.wout(w53_25));
	PE pe53_26(.x(x26),.w(w53_25),.acc(r53_25),.res(r53_26),.clk(clk),.wout(w53_26));
	PE pe53_27(.x(x27),.w(w53_26),.acc(r53_26),.res(r53_27),.clk(clk),.wout(w53_27));
	PE pe53_28(.x(x28),.w(w53_27),.acc(r53_27),.res(r53_28),.clk(clk),.wout(w53_28));
	PE pe53_29(.x(x29),.w(w53_28),.acc(r53_28),.res(r53_29),.clk(clk),.wout(w53_29));
	PE pe53_30(.x(x30),.w(w53_29),.acc(r53_29),.res(r53_30),.clk(clk),.wout(w53_30));
	PE pe53_31(.x(x31),.w(w53_30),.acc(r53_30),.res(r53_31),.clk(clk),.wout(w53_31));
	PE pe53_32(.x(x32),.w(w53_31),.acc(r53_31),.res(r53_32),.clk(clk),.wout(w53_32));
	PE pe53_33(.x(x33),.w(w53_32),.acc(r53_32),.res(r53_33),.clk(clk),.wout(w53_33));
	PE pe53_34(.x(x34),.w(w53_33),.acc(r53_33),.res(r53_34),.clk(clk),.wout(w53_34));
	PE pe53_35(.x(x35),.w(w53_34),.acc(r53_34),.res(r53_35),.clk(clk),.wout(w53_35));
	PE pe53_36(.x(x36),.w(w53_35),.acc(r53_35),.res(r53_36),.clk(clk),.wout(w53_36));
	PE pe53_37(.x(x37),.w(w53_36),.acc(r53_36),.res(r53_37),.clk(clk),.wout(w53_37));
	PE pe53_38(.x(x38),.w(w53_37),.acc(r53_37),.res(r53_38),.clk(clk),.wout(w53_38));
	PE pe53_39(.x(x39),.w(w53_38),.acc(r53_38),.res(r53_39),.clk(clk),.wout(w53_39));
	PE pe53_40(.x(x40),.w(w53_39),.acc(r53_39),.res(r53_40),.clk(clk),.wout(w53_40));
	PE pe53_41(.x(x41),.w(w53_40),.acc(r53_40),.res(r53_41),.clk(clk),.wout(w53_41));
	PE pe53_42(.x(x42),.w(w53_41),.acc(r53_41),.res(r53_42),.clk(clk),.wout(w53_42));
	PE pe53_43(.x(x43),.w(w53_42),.acc(r53_42),.res(r53_43),.clk(clk),.wout(w53_43));
	PE pe53_44(.x(x44),.w(w53_43),.acc(r53_43),.res(r53_44),.clk(clk),.wout(w53_44));
	PE pe53_45(.x(x45),.w(w53_44),.acc(r53_44),.res(r53_45),.clk(clk),.wout(w53_45));
	PE pe53_46(.x(x46),.w(w53_45),.acc(r53_45),.res(r53_46),.clk(clk),.wout(w53_46));
	PE pe53_47(.x(x47),.w(w53_46),.acc(r53_46),.res(r53_47),.clk(clk),.wout(w53_47));
	PE pe53_48(.x(x48),.w(w53_47),.acc(r53_47),.res(r53_48),.clk(clk),.wout(w53_48));
	PE pe53_49(.x(x49),.w(w53_48),.acc(r53_48),.res(r53_49),.clk(clk),.wout(w53_49));
	PE pe53_50(.x(x50),.w(w53_49),.acc(r53_49),.res(r53_50),.clk(clk),.wout(w53_50));
	PE pe53_51(.x(x51),.w(w53_50),.acc(r53_50),.res(r53_51),.clk(clk),.wout(w53_51));
	PE pe53_52(.x(x52),.w(w53_51),.acc(r53_51),.res(r53_52),.clk(clk),.wout(w53_52));
	PE pe53_53(.x(x53),.w(w53_52),.acc(r53_52),.res(r53_53),.clk(clk),.wout(w53_53));
	PE pe53_54(.x(x54),.w(w53_53),.acc(r53_53),.res(r53_54),.clk(clk),.wout(w53_54));
	PE pe53_55(.x(x55),.w(w53_54),.acc(r53_54),.res(r53_55),.clk(clk),.wout(w53_55));
	PE pe53_56(.x(x56),.w(w53_55),.acc(r53_55),.res(r53_56),.clk(clk),.wout(w53_56));
	PE pe53_57(.x(x57),.w(w53_56),.acc(r53_56),.res(r53_57),.clk(clk),.wout(w53_57));
	PE pe53_58(.x(x58),.w(w53_57),.acc(r53_57),.res(r53_58),.clk(clk),.wout(w53_58));
	PE pe53_59(.x(x59),.w(w53_58),.acc(r53_58),.res(r53_59),.clk(clk),.wout(w53_59));
	PE pe53_60(.x(x60),.w(w53_59),.acc(r53_59),.res(r53_60),.clk(clk),.wout(w53_60));
	PE pe53_61(.x(x61),.w(w53_60),.acc(r53_60),.res(r53_61),.clk(clk),.wout(w53_61));
	PE pe53_62(.x(x62),.w(w53_61),.acc(r53_61),.res(r53_62),.clk(clk),.wout(w53_62));
	PE pe53_63(.x(x63),.w(w53_62),.acc(r53_62),.res(r53_63),.clk(clk),.wout(w53_63));
	PE pe53_64(.x(x64),.w(w53_63),.acc(r53_63),.res(r53_64),.clk(clk),.wout(w53_64));
	PE pe53_65(.x(x65),.w(w53_64),.acc(r53_64),.res(r53_65),.clk(clk),.wout(w53_65));
	PE pe53_66(.x(x66),.w(w53_65),.acc(r53_65),.res(r53_66),.clk(clk),.wout(w53_66));
	PE pe53_67(.x(x67),.w(w53_66),.acc(r53_66),.res(r53_67),.clk(clk),.wout(w53_67));
	PE pe53_68(.x(x68),.w(w53_67),.acc(r53_67),.res(r53_68),.clk(clk),.wout(w53_68));
	PE pe53_69(.x(x69),.w(w53_68),.acc(r53_68),.res(r53_69),.clk(clk),.wout(w53_69));
	PE pe53_70(.x(x70),.w(w53_69),.acc(r53_69),.res(r53_70),.clk(clk),.wout(w53_70));
	PE pe53_71(.x(x71),.w(w53_70),.acc(r53_70),.res(r53_71),.clk(clk),.wout(w53_71));
	PE pe53_72(.x(x72),.w(w53_71),.acc(r53_71),.res(r53_72),.clk(clk),.wout(w53_72));
	PE pe53_73(.x(x73),.w(w53_72),.acc(r53_72),.res(r53_73),.clk(clk),.wout(w53_73));
	PE pe53_74(.x(x74),.w(w53_73),.acc(r53_73),.res(r53_74),.clk(clk),.wout(w53_74));
	PE pe53_75(.x(x75),.w(w53_74),.acc(r53_74),.res(r53_75),.clk(clk),.wout(w53_75));
	PE pe53_76(.x(x76),.w(w53_75),.acc(r53_75),.res(r53_76),.clk(clk),.wout(w53_76));
	PE pe53_77(.x(x77),.w(w53_76),.acc(r53_76),.res(r53_77),.clk(clk),.wout(w53_77));
	PE pe53_78(.x(x78),.w(w53_77),.acc(r53_77),.res(r53_78),.clk(clk),.wout(w53_78));
	PE pe53_79(.x(x79),.w(w53_78),.acc(r53_78),.res(r53_79),.clk(clk),.wout(w53_79));
	PE pe53_80(.x(x80),.w(w53_79),.acc(r53_79),.res(r53_80),.clk(clk),.wout(w53_80));
	PE pe53_81(.x(x81),.w(w53_80),.acc(r53_80),.res(r53_81),.clk(clk),.wout(w53_81));
	PE pe53_82(.x(x82),.w(w53_81),.acc(r53_81),.res(r53_82),.clk(clk),.wout(w53_82));
	PE pe53_83(.x(x83),.w(w53_82),.acc(r53_82),.res(r53_83),.clk(clk),.wout(w53_83));
	PE pe53_84(.x(x84),.w(w53_83),.acc(r53_83),.res(r53_84),.clk(clk),.wout(w53_84));
	PE pe53_85(.x(x85),.w(w53_84),.acc(r53_84),.res(r53_85),.clk(clk),.wout(w53_85));
	PE pe53_86(.x(x86),.w(w53_85),.acc(r53_85),.res(r53_86),.clk(clk),.wout(w53_86));
	PE pe53_87(.x(x87),.w(w53_86),.acc(r53_86),.res(r53_87),.clk(clk),.wout(w53_87));
	PE pe53_88(.x(x88),.w(w53_87),.acc(r53_87),.res(r53_88),.clk(clk),.wout(w53_88));
	PE pe53_89(.x(x89),.w(w53_88),.acc(r53_88),.res(r53_89),.clk(clk),.wout(w53_89));
	PE pe53_90(.x(x90),.w(w53_89),.acc(r53_89),.res(r53_90),.clk(clk),.wout(w53_90));
	PE pe53_91(.x(x91),.w(w53_90),.acc(r53_90),.res(r53_91),.clk(clk),.wout(w53_91));
	PE pe53_92(.x(x92),.w(w53_91),.acc(r53_91),.res(r53_92),.clk(clk),.wout(w53_92));
	PE pe53_93(.x(x93),.w(w53_92),.acc(r53_92),.res(r53_93),.clk(clk),.wout(w53_93));
	PE pe53_94(.x(x94),.w(w53_93),.acc(r53_93),.res(r53_94),.clk(clk),.wout(w53_94));
	PE pe53_95(.x(x95),.w(w53_94),.acc(r53_94),.res(r53_95),.clk(clk),.wout(w53_95));
	PE pe53_96(.x(x96),.w(w53_95),.acc(r53_95),.res(r53_96),.clk(clk),.wout(w53_96));
	PE pe53_97(.x(x97),.w(w53_96),.acc(r53_96),.res(r53_97),.clk(clk),.wout(w53_97));
	PE pe53_98(.x(x98),.w(w53_97),.acc(r53_97),.res(r53_98),.clk(clk),.wout(w53_98));
	PE pe53_99(.x(x99),.w(w53_98),.acc(r53_98),.res(r53_99),.clk(clk),.wout(w53_99));
	PE pe53_100(.x(x100),.w(w53_99),.acc(r53_99),.res(r53_100),.clk(clk),.wout(w53_100));
	PE pe53_101(.x(x101),.w(w53_100),.acc(r53_100),.res(r53_101),.clk(clk),.wout(w53_101));
	PE pe53_102(.x(x102),.w(w53_101),.acc(r53_101),.res(r53_102),.clk(clk),.wout(w53_102));
	PE pe53_103(.x(x103),.w(w53_102),.acc(r53_102),.res(r53_103),.clk(clk),.wout(w53_103));
	PE pe53_104(.x(x104),.w(w53_103),.acc(r53_103),.res(r53_104),.clk(clk),.wout(w53_104));
	PE pe53_105(.x(x105),.w(w53_104),.acc(r53_104),.res(r53_105),.clk(clk),.wout(w53_105));
	PE pe53_106(.x(x106),.w(w53_105),.acc(r53_105),.res(r53_106),.clk(clk),.wout(w53_106));
	PE pe53_107(.x(x107),.w(w53_106),.acc(r53_106),.res(r53_107),.clk(clk),.wout(w53_107));
	PE pe53_108(.x(x108),.w(w53_107),.acc(r53_107),.res(r53_108),.clk(clk),.wout(w53_108));
	PE pe53_109(.x(x109),.w(w53_108),.acc(r53_108),.res(r53_109),.clk(clk),.wout(w53_109));
	PE pe53_110(.x(x110),.w(w53_109),.acc(r53_109),.res(r53_110),.clk(clk),.wout(w53_110));
	PE pe53_111(.x(x111),.w(w53_110),.acc(r53_110),.res(r53_111),.clk(clk),.wout(w53_111));
	PE pe53_112(.x(x112),.w(w53_111),.acc(r53_111),.res(r53_112),.clk(clk),.wout(w53_112));
	PE pe53_113(.x(x113),.w(w53_112),.acc(r53_112),.res(r53_113),.clk(clk),.wout(w53_113));
	PE pe53_114(.x(x114),.w(w53_113),.acc(r53_113),.res(r53_114),.clk(clk),.wout(w53_114));
	PE pe53_115(.x(x115),.w(w53_114),.acc(r53_114),.res(r53_115),.clk(clk),.wout(w53_115));
	PE pe53_116(.x(x116),.w(w53_115),.acc(r53_115),.res(r53_116),.clk(clk),.wout(w53_116));
	PE pe53_117(.x(x117),.w(w53_116),.acc(r53_116),.res(r53_117),.clk(clk),.wout(w53_117));
	PE pe53_118(.x(x118),.w(w53_117),.acc(r53_117),.res(r53_118),.clk(clk),.wout(w53_118));
	PE pe53_119(.x(x119),.w(w53_118),.acc(r53_118),.res(r53_119),.clk(clk),.wout(w53_119));
	PE pe53_120(.x(x120),.w(w53_119),.acc(r53_119),.res(r53_120),.clk(clk),.wout(w53_120));
	PE pe53_121(.x(x121),.w(w53_120),.acc(r53_120),.res(r53_121),.clk(clk),.wout(w53_121));
	PE pe53_122(.x(x122),.w(w53_121),.acc(r53_121),.res(r53_122),.clk(clk),.wout(w53_122));
	PE pe53_123(.x(x123),.w(w53_122),.acc(r53_122),.res(r53_123),.clk(clk),.wout(w53_123));
	PE pe53_124(.x(x124),.w(w53_123),.acc(r53_123),.res(r53_124),.clk(clk),.wout(w53_124));
	PE pe53_125(.x(x125),.w(w53_124),.acc(r53_124),.res(r53_125),.clk(clk),.wout(w53_125));
	PE pe53_126(.x(x126),.w(w53_125),.acc(r53_125),.res(r53_126),.clk(clk),.wout(w53_126));
	PE pe53_127(.x(x127),.w(w53_126),.acc(r53_126),.res(result53),.clk(clk),.wout(weight53));

	PE pe54_0(.x(x0),.w(w54),.acc(32'h0),.res(r54_0),.clk(clk),.wout(w54_0));
	PE pe54_1(.x(x1),.w(w54_0),.acc(r54_0),.res(r54_1),.clk(clk),.wout(w54_1));
	PE pe54_2(.x(x2),.w(w54_1),.acc(r54_1),.res(r54_2),.clk(clk),.wout(w54_2));
	PE pe54_3(.x(x3),.w(w54_2),.acc(r54_2),.res(r54_3),.clk(clk),.wout(w54_3));
	PE pe54_4(.x(x4),.w(w54_3),.acc(r54_3),.res(r54_4),.clk(clk),.wout(w54_4));
	PE pe54_5(.x(x5),.w(w54_4),.acc(r54_4),.res(r54_5),.clk(clk),.wout(w54_5));
	PE pe54_6(.x(x6),.w(w54_5),.acc(r54_5),.res(r54_6),.clk(clk),.wout(w54_6));
	PE pe54_7(.x(x7),.w(w54_6),.acc(r54_6),.res(r54_7),.clk(clk),.wout(w54_7));
	PE pe54_8(.x(x8),.w(w54_7),.acc(r54_7),.res(r54_8),.clk(clk),.wout(w54_8));
	PE pe54_9(.x(x9),.w(w54_8),.acc(r54_8),.res(r54_9),.clk(clk),.wout(w54_9));
	PE pe54_10(.x(x10),.w(w54_9),.acc(r54_9),.res(r54_10),.clk(clk),.wout(w54_10));
	PE pe54_11(.x(x11),.w(w54_10),.acc(r54_10),.res(r54_11),.clk(clk),.wout(w54_11));
	PE pe54_12(.x(x12),.w(w54_11),.acc(r54_11),.res(r54_12),.clk(clk),.wout(w54_12));
	PE pe54_13(.x(x13),.w(w54_12),.acc(r54_12),.res(r54_13),.clk(clk),.wout(w54_13));
	PE pe54_14(.x(x14),.w(w54_13),.acc(r54_13),.res(r54_14),.clk(clk),.wout(w54_14));
	PE pe54_15(.x(x15),.w(w54_14),.acc(r54_14),.res(r54_15),.clk(clk),.wout(w54_15));
	PE pe54_16(.x(x16),.w(w54_15),.acc(r54_15),.res(r54_16),.clk(clk),.wout(w54_16));
	PE pe54_17(.x(x17),.w(w54_16),.acc(r54_16),.res(r54_17),.clk(clk),.wout(w54_17));
	PE pe54_18(.x(x18),.w(w54_17),.acc(r54_17),.res(r54_18),.clk(clk),.wout(w54_18));
	PE pe54_19(.x(x19),.w(w54_18),.acc(r54_18),.res(r54_19),.clk(clk),.wout(w54_19));
	PE pe54_20(.x(x20),.w(w54_19),.acc(r54_19),.res(r54_20),.clk(clk),.wout(w54_20));
	PE pe54_21(.x(x21),.w(w54_20),.acc(r54_20),.res(r54_21),.clk(clk),.wout(w54_21));
	PE pe54_22(.x(x22),.w(w54_21),.acc(r54_21),.res(r54_22),.clk(clk),.wout(w54_22));
	PE pe54_23(.x(x23),.w(w54_22),.acc(r54_22),.res(r54_23),.clk(clk),.wout(w54_23));
	PE pe54_24(.x(x24),.w(w54_23),.acc(r54_23),.res(r54_24),.clk(clk),.wout(w54_24));
	PE pe54_25(.x(x25),.w(w54_24),.acc(r54_24),.res(r54_25),.clk(clk),.wout(w54_25));
	PE pe54_26(.x(x26),.w(w54_25),.acc(r54_25),.res(r54_26),.clk(clk),.wout(w54_26));
	PE pe54_27(.x(x27),.w(w54_26),.acc(r54_26),.res(r54_27),.clk(clk),.wout(w54_27));
	PE pe54_28(.x(x28),.w(w54_27),.acc(r54_27),.res(r54_28),.clk(clk),.wout(w54_28));
	PE pe54_29(.x(x29),.w(w54_28),.acc(r54_28),.res(r54_29),.clk(clk),.wout(w54_29));
	PE pe54_30(.x(x30),.w(w54_29),.acc(r54_29),.res(r54_30),.clk(clk),.wout(w54_30));
	PE pe54_31(.x(x31),.w(w54_30),.acc(r54_30),.res(r54_31),.clk(clk),.wout(w54_31));
	PE pe54_32(.x(x32),.w(w54_31),.acc(r54_31),.res(r54_32),.clk(clk),.wout(w54_32));
	PE pe54_33(.x(x33),.w(w54_32),.acc(r54_32),.res(r54_33),.clk(clk),.wout(w54_33));
	PE pe54_34(.x(x34),.w(w54_33),.acc(r54_33),.res(r54_34),.clk(clk),.wout(w54_34));
	PE pe54_35(.x(x35),.w(w54_34),.acc(r54_34),.res(r54_35),.clk(clk),.wout(w54_35));
	PE pe54_36(.x(x36),.w(w54_35),.acc(r54_35),.res(r54_36),.clk(clk),.wout(w54_36));
	PE pe54_37(.x(x37),.w(w54_36),.acc(r54_36),.res(r54_37),.clk(clk),.wout(w54_37));
	PE pe54_38(.x(x38),.w(w54_37),.acc(r54_37),.res(r54_38),.clk(clk),.wout(w54_38));
	PE pe54_39(.x(x39),.w(w54_38),.acc(r54_38),.res(r54_39),.clk(clk),.wout(w54_39));
	PE pe54_40(.x(x40),.w(w54_39),.acc(r54_39),.res(r54_40),.clk(clk),.wout(w54_40));
	PE pe54_41(.x(x41),.w(w54_40),.acc(r54_40),.res(r54_41),.clk(clk),.wout(w54_41));
	PE pe54_42(.x(x42),.w(w54_41),.acc(r54_41),.res(r54_42),.clk(clk),.wout(w54_42));
	PE pe54_43(.x(x43),.w(w54_42),.acc(r54_42),.res(r54_43),.clk(clk),.wout(w54_43));
	PE pe54_44(.x(x44),.w(w54_43),.acc(r54_43),.res(r54_44),.clk(clk),.wout(w54_44));
	PE pe54_45(.x(x45),.w(w54_44),.acc(r54_44),.res(r54_45),.clk(clk),.wout(w54_45));
	PE pe54_46(.x(x46),.w(w54_45),.acc(r54_45),.res(r54_46),.clk(clk),.wout(w54_46));
	PE pe54_47(.x(x47),.w(w54_46),.acc(r54_46),.res(r54_47),.clk(clk),.wout(w54_47));
	PE pe54_48(.x(x48),.w(w54_47),.acc(r54_47),.res(r54_48),.clk(clk),.wout(w54_48));
	PE pe54_49(.x(x49),.w(w54_48),.acc(r54_48),.res(r54_49),.clk(clk),.wout(w54_49));
	PE pe54_50(.x(x50),.w(w54_49),.acc(r54_49),.res(r54_50),.clk(clk),.wout(w54_50));
	PE pe54_51(.x(x51),.w(w54_50),.acc(r54_50),.res(r54_51),.clk(clk),.wout(w54_51));
	PE pe54_52(.x(x52),.w(w54_51),.acc(r54_51),.res(r54_52),.clk(clk),.wout(w54_52));
	PE pe54_53(.x(x53),.w(w54_52),.acc(r54_52),.res(r54_53),.clk(clk),.wout(w54_53));
	PE pe54_54(.x(x54),.w(w54_53),.acc(r54_53),.res(r54_54),.clk(clk),.wout(w54_54));
	PE pe54_55(.x(x55),.w(w54_54),.acc(r54_54),.res(r54_55),.clk(clk),.wout(w54_55));
	PE pe54_56(.x(x56),.w(w54_55),.acc(r54_55),.res(r54_56),.clk(clk),.wout(w54_56));
	PE pe54_57(.x(x57),.w(w54_56),.acc(r54_56),.res(r54_57),.clk(clk),.wout(w54_57));
	PE pe54_58(.x(x58),.w(w54_57),.acc(r54_57),.res(r54_58),.clk(clk),.wout(w54_58));
	PE pe54_59(.x(x59),.w(w54_58),.acc(r54_58),.res(r54_59),.clk(clk),.wout(w54_59));
	PE pe54_60(.x(x60),.w(w54_59),.acc(r54_59),.res(r54_60),.clk(clk),.wout(w54_60));
	PE pe54_61(.x(x61),.w(w54_60),.acc(r54_60),.res(r54_61),.clk(clk),.wout(w54_61));
	PE pe54_62(.x(x62),.w(w54_61),.acc(r54_61),.res(r54_62),.clk(clk),.wout(w54_62));
	PE pe54_63(.x(x63),.w(w54_62),.acc(r54_62),.res(r54_63),.clk(clk),.wout(w54_63));
	PE pe54_64(.x(x64),.w(w54_63),.acc(r54_63),.res(r54_64),.clk(clk),.wout(w54_64));
	PE pe54_65(.x(x65),.w(w54_64),.acc(r54_64),.res(r54_65),.clk(clk),.wout(w54_65));
	PE pe54_66(.x(x66),.w(w54_65),.acc(r54_65),.res(r54_66),.clk(clk),.wout(w54_66));
	PE pe54_67(.x(x67),.w(w54_66),.acc(r54_66),.res(r54_67),.clk(clk),.wout(w54_67));
	PE pe54_68(.x(x68),.w(w54_67),.acc(r54_67),.res(r54_68),.clk(clk),.wout(w54_68));
	PE pe54_69(.x(x69),.w(w54_68),.acc(r54_68),.res(r54_69),.clk(clk),.wout(w54_69));
	PE pe54_70(.x(x70),.w(w54_69),.acc(r54_69),.res(r54_70),.clk(clk),.wout(w54_70));
	PE pe54_71(.x(x71),.w(w54_70),.acc(r54_70),.res(r54_71),.clk(clk),.wout(w54_71));
	PE pe54_72(.x(x72),.w(w54_71),.acc(r54_71),.res(r54_72),.clk(clk),.wout(w54_72));
	PE pe54_73(.x(x73),.w(w54_72),.acc(r54_72),.res(r54_73),.clk(clk),.wout(w54_73));
	PE pe54_74(.x(x74),.w(w54_73),.acc(r54_73),.res(r54_74),.clk(clk),.wout(w54_74));
	PE pe54_75(.x(x75),.w(w54_74),.acc(r54_74),.res(r54_75),.clk(clk),.wout(w54_75));
	PE pe54_76(.x(x76),.w(w54_75),.acc(r54_75),.res(r54_76),.clk(clk),.wout(w54_76));
	PE pe54_77(.x(x77),.w(w54_76),.acc(r54_76),.res(r54_77),.clk(clk),.wout(w54_77));
	PE pe54_78(.x(x78),.w(w54_77),.acc(r54_77),.res(r54_78),.clk(clk),.wout(w54_78));
	PE pe54_79(.x(x79),.w(w54_78),.acc(r54_78),.res(r54_79),.clk(clk),.wout(w54_79));
	PE pe54_80(.x(x80),.w(w54_79),.acc(r54_79),.res(r54_80),.clk(clk),.wout(w54_80));
	PE pe54_81(.x(x81),.w(w54_80),.acc(r54_80),.res(r54_81),.clk(clk),.wout(w54_81));
	PE pe54_82(.x(x82),.w(w54_81),.acc(r54_81),.res(r54_82),.clk(clk),.wout(w54_82));
	PE pe54_83(.x(x83),.w(w54_82),.acc(r54_82),.res(r54_83),.clk(clk),.wout(w54_83));
	PE pe54_84(.x(x84),.w(w54_83),.acc(r54_83),.res(r54_84),.clk(clk),.wout(w54_84));
	PE pe54_85(.x(x85),.w(w54_84),.acc(r54_84),.res(r54_85),.clk(clk),.wout(w54_85));
	PE pe54_86(.x(x86),.w(w54_85),.acc(r54_85),.res(r54_86),.clk(clk),.wout(w54_86));
	PE pe54_87(.x(x87),.w(w54_86),.acc(r54_86),.res(r54_87),.clk(clk),.wout(w54_87));
	PE pe54_88(.x(x88),.w(w54_87),.acc(r54_87),.res(r54_88),.clk(clk),.wout(w54_88));
	PE pe54_89(.x(x89),.w(w54_88),.acc(r54_88),.res(r54_89),.clk(clk),.wout(w54_89));
	PE pe54_90(.x(x90),.w(w54_89),.acc(r54_89),.res(r54_90),.clk(clk),.wout(w54_90));
	PE pe54_91(.x(x91),.w(w54_90),.acc(r54_90),.res(r54_91),.clk(clk),.wout(w54_91));
	PE pe54_92(.x(x92),.w(w54_91),.acc(r54_91),.res(r54_92),.clk(clk),.wout(w54_92));
	PE pe54_93(.x(x93),.w(w54_92),.acc(r54_92),.res(r54_93),.clk(clk),.wout(w54_93));
	PE pe54_94(.x(x94),.w(w54_93),.acc(r54_93),.res(r54_94),.clk(clk),.wout(w54_94));
	PE pe54_95(.x(x95),.w(w54_94),.acc(r54_94),.res(r54_95),.clk(clk),.wout(w54_95));
	PE pe54_96(.x(x96),.w(w54_95),.acc(r54_95),.res(r54_96),.clk(clk),.wout(w54_96));
	PE pe54_97(.x(x97),.w(w54_96),.acc(r54_96),.res(r54_97),.clk(clk),.wout(w54_97));
	PE pe54_98(.x(x98),.w(w54_97),.acc(r54_97),.res(r54_98),.clk(clk),.wout(w54_98));
	PE pe54_99(.x(x99),.w(w54_98),.acc(r54_98),.res(r54_99),.clk(clk),.wout(w54_99));
	PE pe54_100(.x(x100),.w(w54_99),.acc(r54_99),.res(r54_100),.clk(clk),.wout(w54_100));
	PE pe54_101(.x(x101),.w(w54_100),.acc(r54_100),.res(r54_101),.clk(clk),.wout(w54_101));
	PE pe54_102(.x(x102),.w(w54_101),.acc(r54_101),.res(r54_102),.clk(clk),.wout(w54_102));
	PE pe54_103(.x(x103),.w(w54_102),.acc(r54_102),.res(r54_103),.clk(clk),.wout(w54_103));
	PE pe54_104(.x(x104),.w(w54_103),.acc(r54_103),.res(r54_104),.clk(clk),.wout(w54_104));
	PE pe54_105(.x(x105),.w(w54_104),.acc(r54_104),.res(r54_105),.clk(clk),.wout(w54_105));
	PE pe54_106(.x(x106),.w(w54_105),.acc(r54_105),.res(r54_106),.clk(clk),.wout(w54_106));
	PE pe54_107(.x(x107),.w(w54_106),.acc(r54_106),.res(r54_107),.clk(clk),.wout(w54_107));
	PE pe54_108(.x(x108),.w(w54_107),.acc(r54_107),.res(r54_108),.clk(clk),.wout(w54_108));
	PE pe54_109(.x(x109),.w(w54_108),.acc(r54_108),.res(r54_109),.clk(clk),.wout(w54_109));
	PE pe54_110(.x(x110),.w(w54_109),.acc(r54_109),.res(r54_110),.clk(clk),.wout(w54_110));
	PE pe54_111(.x(x111),.w(w54_110),.acc(r54_110),.res(r54_111),.clk(clk),.wout(w54_111));
	PE pe54_112(.x(x112),.w(w54_111),.acc(r54_111),.res(r54_112),.clk(clk),.wout(w54_112));
	PE pe54_113(.x(x113),.w(w54_112),.acc(r54_112),.res(r54_113),.clk(clk),.wout(w54_113));
	PE pe54_114(.x(x114),.w(w54_113),.acc(r54_113),.res(r54_114),.clk(clk),.wout(w54_114));
	PE pe54_115(.x(x115),.w(w54_114),.acc(r54_114),.res(r54_115),.clk(clk),.wout(w54_115));
	PE pe54_116(.x(x116),.w(w54_115),.acc(r54_115),.res(r54_116),.clk(clk),.wout(w54_116));
	PE pe54_117(.x(x117),.w(w54_116),.acc(r54_116),.res(r54_117),.clk(clk),.wout(w54_117));
	PE pe54_118(.x(x118),.w(w54_117),.acc(r54_117),.res(r54_118),.clk(clk),.wout(w54_118));
	PE pe54_119(.x(x119),.w(w54_118),.acc(r54_118),.res(r54_119),.clk(clk),.wout(w54_119));
	PE pe54_120(.x(x120),.w(w54_119),.acc(r54_119),.res(r54_120),.clk(clk),.wout(w54_120));
	PE pe54_121(.x(x121),.w(w54_120),.acc(r54_120),.res(r54_121),.clk(clk),.wout(w54_121));
	PE pe54_122(.x(x122),.w(w54_121),.acc(r54_121),.res(r54_122),.clk(clk),.wout(w54_122));
	PE pe54_123(.x(x123),.w(w54_122),.acc(r54_122),.res(r54_123),.clk(clk),.wout(w54_123));
	PE pe54_124(.x(x124),.w(w54_123),.acc(r54_123),.res(r54_124),.clk(clk),.wout(w54_124));
	PE pe54_125(.x(x125),.w(w54_124),.acc(r54_124),.res(r54_125),.clk(clk),.wout(w54_125));
	PE pe54_126(.x(x126),.w(w54_125),.acc(r54_125),.res(r54_126),.clk(clk),.wout(w54_126));
	PE pe54_127(.x(x127),.w(w54_126),.acc(r54_126),.res(result54),.clk(clk),.wout(weight54));

	PE pe55_0(.x(x0),.w(w55),.acc(32'h0),.res(r55_0),.clk(clk),.wout(w55_0));
	PE pe55_1(.x(x1),.w(w55_0),.acc(r55_0),.res(r55_1),.clk(clk),.wout(w55_1));
	PE pe55_2(.x(x2),.w(w55_1),.acc(r55_1),.res(r55_2),.clk(clk),.wout(w55_2));
	PE pe55_3(.x(x3),.w(w55_2),.acc(r55_2),.res(r55_3),.clk(clk),.wout(w55_3));
	PE pe55_4(.x(x4),.w(w55_3),.acc(r55_3),.res(r55_4),.clk(clk),.wout(w55_4));
	PE pe55_5(.x(x5),.w(w55_4),.acc(r55_4),.res(r55_5),.clk(clk),.wout(w55_5));
	PE pe55_6(.x(x6),.w(w55_5),.acc(r55_5),.res(r55_6),.clk(clk),.wout(w55_6));
	PE pe55_7(.x(x7),.w(w55_6),.acc(r55_6),.res(r55_7),.clk(clk),.wout(w55_7));
	PE pe55_8(.x(x8),.w(w55_7),.acc(r55_7),.res(r55_8),.clk(clk),.wout(w55_8));
	PE pe55_9(.x(x9),.w(w55_8),.acc(r55_8),.res(r55_9),.clk(clk),.wout(w55_9));
	PE pe55_10(.x(x10),.w(w55_9),.acc(r55_9),.res(r55_10),.clk(clk),.wout(w55_10));
	PE pe55_11(.x(x11),.w(w55_10),.acc(r55_10),.res(r55_11),.clk(clk),.wout(w55_11));
	PE pe55_12(.x(x12),.w(w55_11),.acc(r55_11),.res(r55_12),.clk(clk),.wout(w55_12));
	PE pe55_13(.x(x13),.w(w55_12),.acc(r55_12),.res(r55_13),.clk(clk),.wout(w55_13));
	PE pe55_14(.x(x14),.w(w55_13),.acc(r55_13),.res(r55_14),.clk(clk),.wout(w55_14));
	PE pe55_15(.x(x15),.w(w55_14),.acc(r55_14),.res(r55_15),.clk(clk),.wout(w55_15));
	PE pe55_16(.x(x16),.w(w55_15),.acc(r55_15),.res(r55_16),.clk(clk),.wout(w55_16));
	PE pe55_17(.x(x17),.w(w55_16),.acc(r55_16),.res(r55_17),.clk(clk),.wout(w55_17));
	PE pe55_18(.x(x18),.w(w55_17),.acc(r55_17),.res(r55_18),.clk(clk),.wout(w55_18));
	PE pe55_19(.x(x19),.w(w55_18),.acc(r55_18),.res(r55_19),.clk(clk),.wout(w55_19));
	PE pe55_20(.x(x20),.w(w55_19),.acc(r55_19),.res(r55_20),.clk(clk),.wout(w55_20));
	PE pe55_21(.x(x21),.w(w55_20),.acc(r55_20),.res(r55_21),.clk(clk),.wout(w55_21));
	PE pe55_22(.x(x22),.w(w55_21),.acc(r55_21),.res(r55_22),.clk(clk),.wout(w55_22));
	PE pe55_23(.x(x23),.w(w55_22),.acc(r55_22),.res(r55_23),.clk(clk),.wout(w55_23));
	PE pe55_24(.x(x24),.w(w55_23),.acc(r55_23),.res(r55_24),.clk(clk),.wout(w55_24));
	PE pe55_25(.x(x25),.w(w55_24),.acc(r55_24),.res(r55_25),.clk(clk),.wout(w55_25));
	PE pe55_26(.x(x26),.w(w55_25),.acc(r55_25),.res(r55_26),.clk(clk),.wout(w55_26));
	PE pe55_27(.x(x27),.w(w55_26),.acc(r55_26),.res(r55_27),.clk(clk),.wout(w55_27));
	PE pe55_28(.x(x28),.w(w55_27),.acc(r55_27),.res(r55_28),.clk(clk),.wout(w55_28));
	PE pe55_29(.x(x29),.w(w55_28),.acc(r55_28),.res(r55_29),.clk(clk),.wout(w55_29));
	PE pe55_30(.x(x30),.w(w55_29),.acc(r55_29),.res(r55_30),.clk(clk),.wout(w55_30));
	PE pe55_31(.x(x31),.w(w55_30),.acc(r55_30),.res(r55_31),.clk(clk),.wout(w55_31));
	PE pe55_32(.x(x32),.w(w55_31),.acc(r55_31),.res(r55_32),.clk(clk),.wout(w55_32));
	PE pe55_33(.x(x33),.w(w55_32),.acc(r55_32),.res(r55_33),.clk(clk),.wout(w55_33));
	PE pe55_34(.x(x34),.w(w55_33),.acc(r55_33),.res(r55_34),.clk(clk),.wout(w55_34));
	PE pe55_35(.x(x35),.w(w55_34),.acc(r55_34),.res(r55_35),.clk(clk),.wout(w55_35));
	PE pe55_36(.x(x36),.w(w55_35),.acc(r55_35),.res(r55_36),.clk(clk),.wout(w55_36));
	PE pe55_37(.x(x37),.w(w55_36),.acc(r55_36),.res(r55_37),.clk(clk),.wout(w55_37));
	PE pe55_38(.x(x38),.w(w55_37),.acc(r55_37),.res(r55_38),.clk(clk),.wout(w55_38));
	PE pe55_39(.x(x39),.w(w55_38),.acc(r55_38),.res(r55_39),.clk(clk),.wout(w55_39));
	PE pe55_40(.x(x40),.w(w55_39),.acc(r55_39),.res(r55_40),.clk(clk),.wout(w55_40));
	PE pe55_41(.x(x41),.w(w55_40),.acc(r55_40),.res(r55_41),.clk(clk),.wout(w55_41));
	PE pe55_42(.x(x42),.w(w55_41),.acc(r55_41),.res(r55_42),.clk(clk),.wout(w55_42));
	PE pe55_43(.x(x43),.w(w55_42),.acc(r55_42),.res(r55_43),.clk(clk),.wout(w55_43));
	PE pe55_44(.x(x44),.w(w55_43),.acc(r55_43),.res(r55_44),.clk(clk),.wout(w55_44));
	PE pe55_45(.x(x45),.w(w55_44),.acc(r55_44),.res(r55_45),.clk(clk),.wout(w55_45));
	PE pe55_46(.x(x46),.w(w55_45),.acc(r55_45),.res(r55_46),.clk(clk),.wout(w55_46));
	PE pe55_47(.x(x47),.w(w55_46),.acc(r55_46),.res(r55_47),.clk(clk),.wout(w55_47));
	PE pe55_48(.x(x48),.w(w55_47),.acc(r55_47),.res(r55_48),.clk(clk),.wout(w55_48));
	PE pe55_49(.x(x49),.w(w55_48),.acc(r55_48),.res(r55_49),.clk(clk),.wout(w55_49));
	PE pe55_50(.x(x50),.w(w55_49),.acc(r55_49),.res(r55_50),.clk(clk),.wout(w55_50));
	PE pe55_51(.x(x51),.w(w55_50),.acc(r55_50),.res(r55_51),.clk(clk),.wout(w55_51));
	PE pe55_52(.x(x52),.w(w55_51),.acc(r55_51),.res(r55_52),.clk(clk),.wout(w55_52));
	PE pe55_53(.x(x53),.w(w55_52),.acc(r55_52),.res(r55_53),.clk(clk),.wout(w55_53));
	PE pe55_54(.x(x54),.w(w55_53),.acc(r55_53),.res(r55_54),.clk(clk),.wout(w55_54));
	PE pe55_55(.x(x55),.w(w55_54),.acc(r55_54),.res(r55_55),.clk(clk),.wout(w55_55));
	PE pe55_56(.x(x56),.w(w55_55),.acc(r55_55),.res(r55_56),.clk(clk),.wout(w55_56));
	PE pe55_57(.x(x57),.w(w55_56),.acc(r55_56),.res(r55_57),.clk(clk),.wout(w55_57));
	PE pe55_58(.x(x58),.w(w55_57),.acc(r55_57),.res(r55_58),.clk(clk),.wout(w55_58));
	PE pe55_59(.x(x59),.w(w55_58),.acc(r55_58),.res(r55_59),.clk(clk),.wout(w55_59));
	PE pe55_60(.x(x60),.w(w55_59),.acc(r55_59),.res(r55_60),.clk(clk),.wout(w55_60));
	PE pe55_61(.x(x61),.w(w55_60),.acc(r55_60),.res(r55_61),.clk(clk),.wout(w55_61));
	PE pe55_62(.x(x62),.w(w55_61),.acc(r55_61),.res(r55_62),.clk(clk),.wout(w55_62));
	PE pe55_63(.x(x63),.w(w55_62),.acc(r55_62),.res(r55_63),.clk(clk),.wout(w55_63));
	PE pe55_64(.x(x64),.w(w55_63),.acc(r55_63),.res(r55_64),.clk(clk),.wout(w55_64));
	PE pe55_65(.x(x65),.w(w55_64),.acc(r55_64),.res(r55_65),.clk(clk),.wout(w55_65));
	PE pe55_66(.x(x66),.w(w55_65),.acc(r55_65),.res(r55_66),.clk(clk),.wout(w55_66));
	PE pe55_67(.x(x67),.w(w55_66),.acc(r55_66),.res(r55_67),.clk(clk),.wout(w55_67));
	PE pe55_68(.x(x68),.w(w55_67),.acc(r55_67),.res(r55_68),.clk(clk),.wout(w55_68));
	PE pe55_69(.x(x69),.w(w55_68),.acc(r55_68),.res(r55_69),.clk(clk),.wout(w55_69));
	PE pe55_70(.x(x70),.w(w55_69),.acc(r55_69),.res(r55_70),.clk(clk),.wout(w55_70));
	PE pe55_71(.x(x71),.w(w55_70),.acc(r55_70),.res(r55_71),.clk(clk),.wout(w55_71));
	PE pe55_72(.x(x72),.w(w55_71),.acc(r55_71),.res(r55_72),.clk(clk),.wout(w55_72));
	PE pe55_73(.x(x73),.w(w55_72),.acc(r55_72),.res(r55_73),.clk(clk),.wout(w55_73));
	PE pe55_74(.x(x74),.w(w55_73),.acc(r55_73),.res(r55_74),.clk(clk),.wout(w55_74));
	PE pe55_75(.x(x75),.w(w55_74),.acc(r55_74),.res(r55_75),.clk(clk),.wout(w55_75));
	PE pe55_76(.x(x76),.w(w55_75),.acc(r55_75),.res(r55_76),.clk(clk),.wout(w55_76));
	PE pe55_77(.x(x77),.w(w55_76),.acc(r55_76),.res(r55_77),.clk(clk),.wout(w55_77));
	PE pe55_78(.x(x78),.w(w55_77),.acc(r55_77),.res(r55_78),.clk(clk),.wout(w55_78));
	PE pe55_79(.x(x79),.w(w55_78),.acc(r55_78),.res(r55_79),.clk(clk),.wout(w55_79));
	PE pe55_80(.x(x80),.w(w55_79),.acc(r55_79),.res(r55_80),.clk(clk),.wout(w55_80));
	PE pe55_81(.x(x81),.w(w55_80),.acc(r55_80),.res(r55_81),.clk(clk),.wout(w55_81));
	PE pe55_82(.x(x82),.w(w55_81),.acc(r55_81),.res(r55_82),.clk(clk),.wout(w55_82));
	PE pe55_83(.x(x83),.w(w55_82),.acc(r55_82),.res(r55_83),.clk(clk),.wout(w55_83));
	PE pe55_84(.x(x84),.w(w55_83),.acc(r55_83),.res(r55_84),.clk(clk),.wout(w55_84));
	PE pe55_85(.x(x85),.w(w55_84),.acc(r55_84),.res(r55_85),.clk(clk),.wout(w55_85));
	PE pe55_86(.x(x86),.w(w55_85),.acc(r55_85),.res(r55_86),.clk(clk),.wout(w55_86));
	PE pe55_87(.x(x87),.w(w55_86),.acc(r55_86),.res(r55_87),.clk(clk),.wout(w55_87));
	PE pe55_88(.x(x88),.w(w55_87),.acc(r55_87),.res(r55_88),.clk(clk),.wout(w55_88));
	PE pe55_89(.x(x89),.w(w55_88),.acc(r55_88),.res(r55_89),.clk(clk),.wout(w55_89));
	PE pe55_90(.x(x90),.w(w55_89),.acc(r55_89),.res(r55_90),.clk(clk),.wout(w55_90));
	PE pe55_91(.x(x91),.w(w55_90),.acc(r55_90),.res(r55_91),.clk(clk),.wout(w55_91));
	PE pe55_92(.x(x92),.w(w55_91),.acc(r55_91),.res(r55_92),.clk(clk),.wout(w55_92));
	PE pe55_93(.x(x93),.w(w55_92),.acc(r55_92),.res(r55_93),.clk(clk),.wout(w55_93));
	PE pe55_94(.x(x94),.w(w55_93),.acc(r55_93),.res(r55_94),.clk(clk),.wout(w55_94));
	PE pe55_95(.x(x95),.w(w55_94),.acc(r55_94),.res(r55_95),.clk(clk),.wout(w55_95));
	PE pe55_96(.x(x96),.w(w55_95),.acc(r55_95),.res(r55_96),.clk(clk),.wout(w55_96));
	PE pe55_97(.x(x97),.w(w55_96),.acc(r55_96),.res(r55_97),.clk(clk),.wout(w55_97));
	PE pe55_98(.x(x98),.w(w55_97),.acc(r55_97),.res(r55_98),.clk(clk),.wout(w55_98));
	PE pe55_99(.x(x99),.w(w55_98),.acc(r55_98),.res(r55_99),.clk(clk),.wout(w55_99));
	PE pe55_100(.x(x100),.w(w55_99),.acc(r55_99),.res(r55_100),.clk(clk),.wout(w55_100));
	PE pe55_101(.x(x101),.w(w55_100),.acc(r55_100),.res(r55_101),.clk(clk),.wout(w55_101));
	PE pe55_102(.x(x102),.w(w55_101),.acc(r55_101),.res(r55_102),.clk(clk),.wout(w55_102));
	PE pe55_103(.x(x103),.w(w55_102),.acc(r55_102),.res(r55_103),.clk(clk),.wout(w55_103));
	PE pe55_104(.x(x104),.w(w55_103),.acc(r55_103),.res(r55_104),.clk(clk),.wout(w55_104));
	PE pe55_105(.x(x105),.w(w55_104),.acc(r55_104),.res(r55_105),.clk(clk),.wout(w55_105));
	PE pe55_106(.x(x106),.w(w55_105),.acc(r55_105),.res(r55_106),.clk(clk),.wout(w55_106));
	PE pe55_107(.x(x107),.w(w55_106),.acc(r55_106),.res(r55_107),.clk(clk),.wout(w55_107));
	PE pe55_108(.x(x108),.w(w55_107),.acc(r55_107),.res(r55_108),.clk(clk),.wout(w55_108));
	PE pe55_109(.x(x109),.w(w55_108),.acc(r55_108),.res(r55_109),.clk(clk),.wout(w55_109));
	PE pe55_110(.x(x110),.w(w55_109),.acc(r55_109),.res(r55_110),.clk(clk),.wout(w55_110));
	PE pe55_111(.x(x111),.w(w55_110),.acc(r55_110),.res(r55_111),.clk(clk),.wout(w55_111));
	PE pe55_112(.x(x112),.w(w55_111),.acc(r55_111),.res(r55_112),.clk(clk),.wout(w55_112));
	PE pe55_113(.x(x113),.w(w55_112),.acc(r55_112),.res(r55_113),.clk(clk),.wout(w55_113));
	PE pe55_114(.x(x114),.w(w55_113),.acc(r55_113),.res(r55_114),.clk(clk),.wout(w55_114));
	PE pe55_115(.x(x115),.w(w55_114),.acc(r55_114),.res(r55_115),.clk(clk),.wout(w55_115));
	PE pe55_116(.x(x116),.w(w55_115),.acc(r55_115),.res(r55_116),.clk(clk),.wout(w55_116));
	PE pe55_117(.x(x117),.w(w55_116),.acc(r55_116),.res(r55_117),.clk(clk),.wout(w55_117));
	PE pe55_118(.x(x118),.w(w55_117),.acc(r55_117),.res(r55_118),.clk(clk),.wout(w55_118));
	PE pe55_119(.x(x119),.w(w55_118),.acc(r55_118),.res(r55_119),.clk(clk),.wout(w55_119));
	PE pe55_120(.x(x120),.w(w55_119),.acc(r55_119),.res(r55_120),.clk(clk),.wout(w55_120));
	PE pe55_121(.x(x121),.w(w55_120),.acc(r55_120),.res(r55_121),.clk(clk),.wout(w55_121));
	PE pe55_122(.x(x122),.w(w55_121),.acc(r55_121),.res(r55_122),.clk(clk),.wout(w55_122));
	PE pe55_123(.x(x123),.w(w55_122),.acc(r55_122),.res(r55_123),.clk(clk),.wout(w55_123));
	PE pe55_124(.x(x124),.w(w55_123),.acc(r55_123),.res(r55_124),.clk(clk),.wout(w55_124));
	PE pe55_125(.x(x125),.w(w55_124),.acc(r55_124),.res(r55_125),.clk(clk),.wout(w55_125));
	PE pe55_126(.x(x126),.w(w55_125),.acc(r55_125),.res(r55_126),.clk(clk),.wout(w55_126));
	PE pe55_127(.x(x127),.w(w55_126),.acc(r55_126),.res(result55),.clk(clk),.wout(weight55));

	PE pe56_0(.x(x0),.w(w56),.acc(32'h0),.res(r56_0),.clk(clk),.wout(w56_0));
	PE pe56_1(.x(x1),.w(w56_0),.acc(r56_0),.res(r56_1),.clk(clk),.wout(w56_1));
	PE pe56_2(.x(x2),.w(w56_1),.acc(r56_1),.res(r56_2),.clk(clk),.wout(w56_2));
	PE pe56_3(.x(x3),.w(w56_2),.acc(r56_2),.res(r56_3),.clk(clk),.wout(w56_3));
	PE pe56_4(.x(x4),.w(w56_3),.acc(r56_3),.res(r56_4),.clk(clk),.wout(w56_4));
	PE pe56_5(.x(x5),.w(w56_4),.acc(r56_4),.res(r56_5),.clk(clk),.wout(w56_5));
	PE pe56_6(.x(x6),.w(w56_5),.acc(r56_5),.res(r56_6),.clk(clk),.wout(w56_6));
	PE pe56_7(.x(x7),.w(w56_6),.acc(r56_6),.res(r56_7),.clk(clk),.wout(w56_7));
	PE pe56_8(.x(x8),.w(w56_7),.acc(r56_7),.res(r56_8),.clk(clk),.wout(w56_8));
	PE pe56_9(.x(x9),.w(w56_8),.acc(r56_8),.res(r56_9),.clk(clk),.wout(w56_9));
	PE pe56_10(.x(x10),.w(w56_9),.acc(r56_9),.res(r56_10),.clk(clk),.wout(w56_10));
	PE pe56_11(.x(x11),.w(w56_10),.acc(r56_10),.res(r56_11),.clk(clk),.wout(w56_11));
	PE pe56_12(.x(x12),.w(w56_11),.acc(r56_11),.res(r56_12),.clk(clk),.wout(w56_12));
	PE pe56_13(.x(x13),.w(w56_12),.acc(r56_12),.res(r56_13),.clk(clk),.wout(w56_13));
	PE pe56_14(.x(x14),.w(w56_13),.acc(r56_13),.res(r56_14),.clk(clk),.wout(w56_14));
	PE pe56_15(.x(x15),.w(w56_14),.acc(r56_14),.res(r56_15),.clk(clk),.wout(w56_15));
	PE pe56_16(.x(x16),.w(w56_15),.acc(r56_15),.res(r56_16),.clk(clk),.wout(w56_16));
	PE pe56_17(.x(x17),.w(w56_16),.acc(r56_16),.res(r56_17),.clk(clk),.wout(w56_17));
	PE pe56_18(.x(x18),.w(w56_17),.acc(r56_17),.res(r56_18),.clk(clk),.wout(w56_18));
	PE pe56_19(.x(x19),.w(w56_18),.acc(r56_18),.res(r56_19),.clk(clk),.wout(w56_19));
	PE pe56_20(.x(x20),.w(w56_19),.acc(r56_19),.res(r56_20),.clk(clk),.wout(w56_20));
	PE pe56_21(.x(x21),.w(w56_20),.acc(r56_20),.res(r56_21),.clk(clk),.wout(w56_21));
	PE pe56_22(.x(x22),.w(w56_21),.acc(r56_21),.res(r56_22),.clk(clk),.wout(w56_22));
	PE pe56_23(.x(x23),.w(w56_22),.acc(r56_22),.res(r56_23),.clk(clk),.wout(w56_23));
	PE pe56_24(.x(x24),.w(w56_23),.acc(r56_23),.res(r56_24),.clk(clk),.wout(w56_24));
	PE pe56_25(.x(x25),.w(w56_24),.acc(r56_24),.res(r56_25),.clk(clk),.wout(w56_25));
	PE pe56_26(.x(x26),.w(w56_25),.acc(r56_25),.res(r56_26),.clk(clk),.wout(w56_26));
	PE pe56_27(.x(x27),.w(w56_26),.acc(r56_26),.res(r56_27),.clk(clk),.wout(w56_27));
	PE pe56_28(.x(x28),.w(w56_27),.acc(r56_27),.res(r56_28),.clk(clk),.wout(w56_28));
	PE pe56_29(.x(x29),.w(w56_28),.acc(r56_28),.res(r56_29),.clk(clk),.wout(w56_29));
	PE pe56_30(.x(x30),.w(w56_29),.acc(r56_29),.res(r56_30),.clk(clk),.wout(w56_30));
	PE pe56_31(.x(x31),.w(w56_30),.acc(r56_30),.res(r56_31),.clk(clk),.wout(w56_31));
	PE pe56_32(.x(x32),.w(w56_31),.acc(r56_31),.res(r56_32),.clk(clk),.wout(w56_32));
	PE pe56_33(.x(x33),.w(w56_32),.acc(r56_32),.res(r56_33),.clk(clk),.wout(w56_33));
	PE pe56_34(.x(x34),.w(w56_33),.acc(r56_33),.res(r56_34),.clk(clk),.wout(w56_34));
	PE pe56_35(.x(x35),.w(w56_34),.acc(r56_34),.res(r56_35),.clk(clk),.wout(w56_35));
	PE pe56_36(.x(x36),.w(w56_35),.acc(r56_35),.res(r56_36),.clk(clk),.wout(w56_36));
	PE pe56_37(.x(x37),.w(w56_36),.acc(r56_36),.res(r56_37),.clk(clk),.wout(w56_37));
	PE pe56_38(.x(x38),.w(w56_37),.acc(r56_37),.res(r56_38),.clk(clk),.wout(w56_38));
	PE pe56_39(.x(x39),.w(w56_38),.acc(r56_38),.res(r56_39),.clk(clk),.wout(w56_39));
	PE pe56_40(.x(x40),.w(w56_39),.acc(r56_39),.res(r56_40),.clk(clk),.wout(w56_40));
	PE pe56_41(.x(x41),.w(w56_40),.acc(r56_40),.res(r56_41),.clk(clk),.wout(w56_41));
	PE pe56_42(.x(x42),.w(w56_41),.acc(r56_41),.res(r56_42),.clk(clk),.wout(w56_42));
	PE pe56_43(.x(x43),.w(w56_42),.acc(r56_42),.res(r56_43),.clk(clk),.wout(w56_43));
	PE pe56_44(.x(x44),.w(w56_43),.acc(r56_43),.res(r56_44),.clk(clk),.wout(w56_44));
	PE pe56_45(.x(x45),.w(w56_44),.acc(r56_44),.res(r56_45),.clk(clk),.wout(w56_45));
	PE pe56_46(.x(x46),.w(w56_45),.acc(r56_45),.res(r56_46),.clk(clk),.wout(w56_46));
	PE pe56_47(.x(x47),.w(w56_46),.acc(r56_46),.res(r56_47),.clk(clk),.wout(w56_47));
	PE pe56_48(.x(x48),.w(w56_47),.acc(r56_47),.res(r56_48),.clk(clk),.wout(w56_48));
	PE pe56_49(.x(x49),.w(w56_48),.acc(r56_48),.res(r56_49),.clk(clk),.wout(w56_49));
	PE pe56_50(.x(x50),.w(w56_49),.acc(r56_49),.res(r56_50),.clk(clk),.wout(w56_50));
	PE pe56_51(.x(x51),.w(w56_50),.acc(r56_50),.res(r56_51),.clk(clk),.wout(w56_51));
	PE pe56_52(.x(x52),.w(w56_51),.acc(r56_51),.res(r56_52),.clk(clk),.wout(w56_52));
	PE pe56_53(.x(x53),.w(w56_52),.acc(r56_52),.res(r56_53),.clk(clk),.wout(w56_53));
	PE pe56_54(.x(x54),.w(w56_53),.acc(r56_53),.res(r56_54),.clk(clk),.wout(w56_54));
	PE pe56_55(.x(x55),.w(w56_54),.acc(r56_54),.res(r56_55),.clk(clk),.wout(w56_55));
	PE pe56_56(.x(x56),.w(w56_55),.acc(r56_55),.res(r56_56),.clk(clk),.wout(w56_56));
	PE pe56_57(.x(x57),.w(w56_56),.acc(r56_56),.res(r56_57),.clk(clk),.wout(w56_57));
	PE pe56_58(.x(x58),.w(w56_57),.acc(r56_57),.res(r56_58),.clk(clk),.wout(w56_58));
	PE pe56_59(.x(x59),.w(w56_58),.acc(r56_58),.res(r56_59),.clk(clk),.wout(w56_59));
	PE pe56_60(.x(x60),.w(w56_59),.acc(r56_59),.res(r56_60),.clk(clk),.wout(w56_60));
	PE pe56_61(.x(x61),.w(w56_60),.acc(r56_60),.res(r56_61),.clk(clk),.wout(w56_61));
	PE pe56_62(.x(x62),.w(w56_61),.acc(r56_61),.res(r56_62),.clk(clk),.wout(w56_62));
	PE pe56_63(.x(x63),.w(w56_62),.acc(r56_62),.res(r56_63),.clk(clk),.wout(w56_63));
	PE pe56_64(.x(x64),.w(w56_63),.acc(r56_63),.res(r56_64),.clk(clk),.wout(w56_64));
	PE pe56_65(.x(x65),.w(w56_64),.acc(r56_64),.res(r56_65),.clk(clk),.wout(w56_65));
	PE pe56_66(.x(x66),.w(w56_65),.acc(r56_65),.res(r56_66),.clk(clk),.wout(w56_66));
	PE pe56_67(.x(x67),.w(w56_66),.acc(r56_66),.res(r56_67),.clk(clk),.wout(w56_67));
	PE pe56_68(.x(x68),.w(w56_67),.acc(r56_67),.res(r56_68),.clk(clk),.wout(w56_68));
	PE pe56_69(.x(x69),.w(w56_68),.acc(r56_68),.res(r56_69),.clk(clk),.wout(w56_69));
	PE pe56_70(.x(x70),.w(w56_69),.acc(r56_69),.res(r56_70),.clk(clk),.wout(w56_70));
	PE pe56_71(.x(x71),.w(w56_70),.acc(r56_70),.res(r56_71),.clk(clk),.wout(w56_71));
	PE pe56_72(.x(x72),.w(w56_71),.acc(r56_71),.res(r56_72),.clk(clk),.wout(w56_72));
	PE pe56_73(.x(x73),.w(w56_72),.acc(r56_72),.res(r56_73),.clk(clk),.wout(w56_73));
	PE pe56_74(.x(x74),.w(w56_73),.acc(r56_73),.res(r56_74),.clk(clk),.wout(w56_74));
	PE pe56_75(.x(x75),.w(w56_74),.acc(r56_74),.res(r56_75),.clk(clk),.wout(w56_75));
	PE pe56_76(.x(x76),.w(w56_75),.acc(r56_75),.res(r56_76),.clk(clk),.wout(w56_76));
	PE pe56_77(.x(x77),.w(w56_76),.acc(r56_76),.res(r56_77),.clk(clk),.wout(w56_77));
	PE pe56_78(.x(x78),.w(w56_77),.acc(r56_77),.res(r56_78),.clk(clk),.wout(w56_78));
	PE pe56_79(.x(x79),.w(w56_78),.acc(r56_78),.res(r56_79),.clk(clk),.wout(w56_79));
	PE pe56_80(.x(x80),.w(w56_79),.acc(r56_79),.res(r56_80),.clk(clk),.wout(w56_80));
	PE pe56_81(.x(x81),.w(w56_80),.acc(r56_80),.res(r56_81),.clk(clk),.wout(w56_81));
	PE pe56_82(.x(x82),.w(w56_81),.acc(r56_81),.res(r56_82),.clk(clk),.wout(w56_82));
	PE pe56_83(.x(x83),.w(w56_82),.acc(r56_82),.res(r56_83),.clk(clk),.wout(w56_83));
	PE pe56_84(.x(x84),.w(w56_83),.acc(r56_83),.res(r56_84),.clk(clk),.wout(w56_84));
	PE pe56_85(.x(x85),.w(w56_84),.acc(r56_84),.res(r56_85),.clk(clk),.wout(w56_85));
	PE pe56_86(.x(x86),.w(w56_85),.acc(r56_85),.res(r56_86),.clk(clk),.wout(w56_86));
	PE pe56_87(.x(x87),.w(w56_86),.acc(r56_86),.res(r56_87),.clk(clk),.wout(w56_87));
	PE pe56_88(.x(x88),.w(w56_87),.acc(r56_87),.res(r56_88),.clk(clk),.wout(w56_88));
	PE pe56_89(.x(x89),.w(w56_88),.acc(r56_88),.res(r56_89),.clk(clk),.wout(w56_89));
	PE pe56_90(.x(x90),.w(w56_89),.acc(r56_89),.res(r56_90),.clk(clk),.wout(w56_90));
	PE pe56_91(.x(x91),.w(w56_90),.acc(r56_90),.res(r56_91),.clk(clk),.wout(w56_91));
	PE pe56_92(.x(x92),.w(w56_91),.acc(r56_91),.res(r56_92),.clk(clk),.wout(w56_92));
	PE pe56_93(.x(x93),.w(w56_92),.acc(r56_92),.res(r56_93),.clk(clk),.wout(w56_93));
	PE pe56_94(.x(x94),.w(w56_93),.acc(r56_93),.res(r56_94),.clk(clk),.wout(w56_94));
	PE pe56_95(.x(x95),.w(w56_94),.acc(r56_94),.res(r56_95),.clk(clk),.wout(w56_95));
	PE pe56_96(.x(x96),.w(w56_95),.acc(r56_95),.res(r56_96),.clk(clk),.wout(w56_96));
	PE pe56_97(.x(x97),.w(w56_96),.acc(r56_96),.res(r56_97),.clk(clk),.wout(w56_97));
	PE pe56_98(.x(x98),.w(w56_97),.acc(r56_97),.res(r56_98),.clk(clk),.wout(w56_98));
	PE pe56_99(.x(x99),.w(w56_98),.acc(r56_98),.res(r56_99),.clk(clk),.wout(w56_99));
	PE pe56_100(.x(x100),.w(w56_99),.acc(r56_99),.res(r56_100),.clk(clk),.wout(w56_100));
	PE pe56_101(.x(x101),.w(w56_100),.acc(r56_100),.res(r56_101),.clk(clk),.wout(w56_101));
	PE pe56_102(.x(x102),.w(w56_101),.acc(r56_101),.res(r56_102),.clk(clk),.wout(w56_102));
	PE pe56_103(.x(x103),.w(w56_102),.acc(r56_102),.res(r56_103),.clk(clk),.wout(w56_103));
	PE pe56_104(.x(x104),.w(w56_103),.acc(r56_103),.res(r56_104),.clk(clk),.wout(w56_104));
	PE pe56_105(.x(x105),.w(w56_104),.acc(r56_104),.res(r56_105),.clk(clk),.wout(w56_105));
	PE pe56_106(.x(x106),.w(w56_105),.acc(r56_105),.res(r56_106),.clk(clk),.wout(w56_106));
	PE pe56_107(.x(x107),.w(w56_106),.acc(r56_106),.res(r56_107),.clk(clk),.wout(w56_107));
	PE pe56_108(.x(x108),.w(w56_107),.acc(r56_107),.res(r56_108),.clk(clk),.wout(w56_108));
	PE pe56_109(.x(x109),.w(w56_108),.acc(r56_108),.res(r56_109),.clk(clk),.wout(w56_109));
	PE pe56_110(.x(x110),.w(w56_109),.acc(r56_109),.res(r56_110),.clk(clk),.wout(w56_110));
	PE pe56_111(.x(x111),.w(w56_110),.acc(r56_110),.res(r56_111),.clk(clk),.wout(w56_111));
	PE pe56_112(.x(x112),.w(w56_111),.acc(r56_111),.res(r56_112),.clk(clk),.wout(w56_112));
	PE pe56_113(.x(x113),.w(w56_112),.acc(r56_112),.res(r56_113),.clk(clk),.wout(w56_113));
	PE pe56_114(.x(x114),.w(w56_113),.acc(r56_113),.res(r56_114),.clk(clk),.wout(w56_114));
	PE pe56_115(.x(x115),.w(w56_114),.acc(r56_114),.res(r56_115),.clk(clk),.wout(w56_115));
	PE pe56_116(.x(x116),.w(w56_115),.acc(r56_115),.res(r56_116),.clk(clk),.wout(w56_116));
	PE pe56_117(.x(x117),.w(w56_116),.acc(r56_116),.res(r56_117),.clk(clk),.wout(w56_117));
	PE pe56_118(.x(x118),.w(w56_117),.acc(r56_117),.res(r56_118),.clk(clk),.wout(w56_118));
	PE pe56_119(.x(x119),.w(w56_118),.acc(r56_118),.res(r56_119),.clk(clk),.wout(w56_119));
	PE pe56_120(.x(x120),.w(w56_119),.acc(r56_119),.res(r56_120),.clk(clk),.wout(w56_120));
	PE pe56_121(.x(x121),.w(w56_120),.acc(r56_120),.res(r56_121),.clk(clk),.wout(w56_121));
	PE pe56_122(.x(x122),.w(w56_121),.acc(r56_121),.res(r56_122),.clk(clk),.wout(w56_122));
	PE pe56_123(.x(x123),.w(w56_122),.acc(r56_122),.res(r56_123),.clk(clk),.wout(w56_123));
	PE pe56_124(.x(x124),.w(w56_123),.acc(r56_123),.res(r56_124),.clk(clk),.wout(w56_124));
	PE pe56_125(.x(x125),.w(w56_124),.acc(r56_124),.res(r56_125),.clk(clk),.wout(w56_125));
	PE pe56_126(.x(x126),.w(w56_125),.acc(r56_125),.res(r56_126),.clk(clk),.wout(w56_126));
	PE pe56_127(.x(x127),.w(w56_126),.acc(r56_126),.res(result56),.clk(clk),.wout(weight56));

	PE pe57_0(.x(x0),.w(w57),.acc(32'h0),.res(r57_0),.clk(clk),.wout(w57_0));
	PE pe57_1(.x(x1),.w(w57_0),.acc(r57_0),.res(r57_1),.clk(clk),.wout(w57_1));
	PE pe57_2(.x(x2),.w(w57_1),.acc(r57_1),.res(r57_2),.clk(clk),.wout(w57_2));
	PE pe57_3(.x(x3),.w(w57_2),.acc(r57_2),.res(r57_3),.clk(clk),.wout(w57_3));
	PE pe57_4(.x(x4),.w(w57_3),.acc(r57_3),.res(r57_4),.clk(clk),.wout(w57_4));
	PE pe57_5(.x(x5),.w(w57_4),.acc(r57_4),.res(r57_5),.clk(clk),.wout(w57_5));
	PE pe57_6(.x(x6),.w(w57_5),.acc(r57_5),.res(r57_6),.clk(clk),.wout(w57_6));
	PE pe57_7(.x(x7),.w(w57_6),.acc(r57_6),.res(r57_7),.clk(clk),.wout(w57_7));
	PE pe57_8(.x(x8),.w(w57_7),.acc(r57_7),.res(r57_8),.clk(clk),.wout(w57_8));
	PE pe57_9(.x(x9),.w(w57_8),.acc(r57_8),.res(r57_9),.clk(clk),.wout(w57_9));
	PE pe57_10(.x(x10),.w(w57_9),.acc(r57_9),.res(r57_10),.clk(clk),.wout(w57_10));
	PE pe57_11(.x(x11),.w(w57_10),.acc(r57_10),.res(r57_11),.clk(clk),.wout(w57_11));
	PE pe57_12(.x(x12),.w(w57_11),.acc(r57_11),.res(r57_12),.clk(clk),.wout(w57_12));
	PE pe57_13(.x(x13),.w(w57_12),.acc(r57_12),.res(r57_13),.clk(clk),.wout(w57_13));
	PE pe57_14(.x(x14),.w(w57_13),.acc(r57_13),.res(r57_14),.clk(clk),.wout(w57_14));
	PE pe57_15(.x(x15),.w(w57_14),.acc(r57_14),.res(r57_15),.clk(clk),.wout(w57_15));
	PE pe57_16(.x(x16),.w(w57_15),.acc(r57_15),.res(r57_16),.clk(clk),.wout(w57_16));
	PE pe57_17(.x(x17),.w(w57_16),.acc(r57_16),.res(r57_17),.clk(clk),.wout(w57_17));
	PE pe57_18(.x(x18),.w(w57_17),.acc(r57_17),.res(r57_18),.clk(clk),.wout(w57_18));
	PE pe57_19(.x(x19),.w(w57_18),.acc(r57_18),.res(r57_19),.clk(clk),.wout(w57_19));
	PE pe57_20(.x(x20),.w(w57_19),.acc(r57_19),.res(r57_20),.clk(clk),.wout(w57_20));
	PE pe57_21(.x(x21),.w(w57_20),.acc(r57_20),.res(r57_21),.clk(clk),.wout(w57_21));
	PE pe57_22(.x(x22),.w(w57_21),.acc(r57_21),.res(r57_22),.clk(clk),.wout(w57_22));
	PE pe57_23(.x(x23),.w(w57_22),.acc(r57_22),.res(r57_23),.clk(clk),.wout(w57_23));
	PE pe57_24(.x(x24),.w(w57_23),.acc(r57_23),.res(r57_24),.clk(clk),.wout(w57_24));
	PE pe57_25(.x(x25),.w(w57_24),.acc(r57_24),.res(r57_25),.clk(clk),.wout(w57_25));
	PE pe57_26(.x(x26),.w(w57_25),.acc(r57_25),.res(r57_26),.clk(clk),.wout(w57_26));
	PE pe57_27(.x(x27),.w(w57_26),.acc(r57_26),.res(r57_27),.clk(clk),.wout(w57_27));
	PE pe57_28(.x(x28),.w(w57_27),.acc(r57_27),.res(r57_28),.clk(clk),.wout(w57_28));
	PE pe57_29(.x(x29),.w(w57_28),.acc(r57_28),.res(r57_29),.clk(clk),.wout(w57_29));
	PE pe57_30(.x(x30),.w(w57_29),.acc(r57_29),.res(r57_30),.clk(clk),.wout(w57_30));
	PE pe57_31(.x(x31),.w(w57_30),.acc(r57_30),.res(r57_31),.clk(clk),.wout(w57_31));
	PE pe57_32(.x(x32),.w(w57_31),.acc(r57_31),.res(r57_32),.clk(clk),.wout(w57_32));
	PE pe57_33(.x(x33),.w(w57_32),.acc(r57_32),.res(r57_33),.clk(clk),.wout(w57_33));
	PE pe57_34(.x(x34),.w(w57_33),.acc(r57_33),.res(r57_34),.clk(clk),.wout(w57_34));
	PE pe57_35(.x(x35),.w(w57_34),.acc(r57_34),.res(r57_35),.clk(clk),.wout(w57_35));
	PE pe57_36(.x(x36),.w(w57_35),.acc(r57_35),.res(r57_36),.clk(clk),.wout(w57_36));
	PE pe57_37(.x(x37),.w(w57_36),.acc(r57_36),.res(r57_37),.clk(clk),.wout(w57_37));
	PE pe57_38(.x(x38),.w(w57_37),.acc(r57_37),.res(r57_38),.clk(clk),.wout(w57_38));
	PE pe57_39(.x(x39),.w(w57_38),.acc(r57_38),.res(r57_39),.clk(clk),.wout(w57_39));
	PE pe57_40(.x(x40),.w(w57_39),.acc(r57_39),.res(r57_40),.clk(clk),.wout(w57_40));
	PE pe57_41(.x(x41),.w(w57_40),.acc(r57_40),.res(r57_41),.clk(clk),.wout(w57_41));
	PE pe57_42(.x(x42),.w(w57_41),.acc(r57_41),.res(r57_42),.clk(clk),.wout(w57_42));
	PE pe57_43(.x(x43),.w(w57_42),.acc(r57_42),.res(r57_43),.clk(clk),.wout(w57_43));
	PE pe57_44(.x(x44),.w(w57_43),.acc(r57_43),.res(r57_44),.clk(clk),.wout(w57_44));
	PE pe57_45(.x(x45),.w(w57_44),.acc(r57_44),.res(r57_45),.clk(clk),.wout(w57_45));
	PE pe57_46(.x(x46),.w(w57_45),.acc(r57_45),.res(r57_46),.clk(clk),.wout(w57_46));
	PE pe57_47(.x(x47),.w(w57_46),.acc(r57_46),.res(r57_47),.clk(clk),.wout(w57_47));
	PE pe57_48(.x(x48),.w(w57_47),.acc(r57_47),.res(r57_48),.clk(clk),.wout(w57_48));
	PE pe57_49(.x(x49),.w(w57_48),.acc(r57_48),.res(r57_49),.clk(clk),.wout(w57_49));
	PE pe57_50(.x(x50),.w(w57_49),.acc(r57_49),.res(r57_50),.clk(clk),.wout(w57_50));
	PE pe57_51(.x(x51),.w(w57_50),.acc(r57_50),.res(r57_51),.clk(clk),.wout(w57_51));
	PE pe57_52(.x(x52),.w(w57_51),.acc(r57_51),.res(r57_52),.clk(clk),.wout(w57_52));
	PE pe57_53(.x(x53),.w(w57_52),.acc(r57_52),.res(r57_53),.clk(clk),.wout(w57_53));
	PE pe57_54(.x(x54),.w(w57_53),.acc(r57_53),.res(r57_54),.clk(clk),.wout(w57_54));
	PE pe57_55(.x(x55),.w(w57_54),.acc(r57_54),.res(r57_55),.clk(clk),.wout(w57_55));
	PE pe57_56(.x(x56),.w(w57_55),.acc(r57_55),.res(r57_56),.clk(clk),.wout(w57_56));
	PE pe57_57(.x(x57),.w(w57_56),.acc(r57_56),.res(r57_57),.clk(clk),.wout(w57_57));
	PE pe57_58(.x(x58),.w(w57_57),.acc(r57_57),.res(r57_58),.clk(clk),.wout(w57_58));
	PE pe57_59(.x(x59),.w(w57_58),.acc(r57_58),.res(r57_59),.clk(clk),.wout(w57_59));
	PE pe57_60(.x(x60),.w(w57_59),.acc(r57_59),.res(r57_60),.clk(clk),.wout(w57_60));
	PE pe57_61(.x(x61),.w(w57_60),.acc(r57_60),.res(r57_61),.clk(clk),.wout(w57_61));
	PE pe57_62(.x(x62),.w(w57_61),.acc(r57_61),.res(r57_62),.clk(clk),.wout(w57_62));
	PE pe57_63(.x(x63),.w(w57_62),.acc(r57_62),.res(r57_63),.clk(clk),.wout(w57_63));
	PE pe57_64(.x(x64),.w(w57_63),.acc(r57_63),.res(r57_64),.clk(clk),.wout(w57_64));
	PE pe57_65(.x(x65),.w(w57_64),.acc(r57_64),.res(r57_65),.clk(clk),.wout(w57_65));
	PE pe57_66(.x(x66),.w(w57_65),.acc(r57_65),.res(r57_66),.clk(clk),.wout(w57_66));
	PE pe57_67(.x(x67),.w(w57_66),.acc(r57_66),.res(r57_67),.clk(clk),.wout(w57_67));
	PE pe57_68(.x(x68),.w(w57_67),.acc(r57_67),.res(r57_68),.clk(clk),.wout(w57_68));
	PE pe57_69(.x(x69),.w(w57_68),.acc(r57_68),.res(r57_69),.clk(clk),.wout(w57_69));
	PE pe57_70(.x(x70),.w(w57_69),.acc(r57_69),.res(r57_70),.clk(clk),.wout(w57_70));
	PE pe57_71(.x(x71),.w(w57_70),.acc(r57_70),.res(r57_71),.clk(clk),.wout(w57_71));
	PE pe57_72(.x(x72),.w(w57_71),.acc(r57_71),.res(r57_72),.clk(clk),.wout(w57_72));
	PE pe57_73(.x(x73),.w(w57_72),.acc(r57_72),.res(r57_73),.clk(clk),.wout(w57_73));
	PE pe57_74(.x(x74),.w(w57_73),.acc(r57_73),.res(r57_74),.clk(clk),.wout(w57_74));
	PE pe57_75(.x(x75),.w(w57_74),.acc(r57_74),.res(r57_75),.clk(clk),.wout(w57_75));
	PE pe57_76(.x(x76),.w(w57_75),.acc(r57_75),.res(r57_76),.clk(clk),.wout(w57_76));
	PE pe57_77(.x(x77),.w(w57_76),.acc(r57_76),.res(r57_77),.clk(clk),.wout(w57_77));
	PE pe57_78(.x(x78),.w(w57_77),.acc(r57_77),.res(r57_78),.clk(clk),.wout(w57_78));
	PE pe57_79(.x(x79),.w(w57_78),.acc(r57_78),.res(r57_79),.clk(clk),.wout(w57_79));
	PE pe57_80(.x(x80),.w(w57_79),.acc(r57_79),.res(r57_80),.clk(clk),.wout(w57_80));
	PE pe57_81(.x(x81),.w(w57_80),.acc(r57_80),.res(r57_81),.clk(clk),.wout(w57_81));
	PE pe57_82(.x(x82),.w(w57_81),.acc(r57_81),.res(r57_82),.clk(clk),.wout(w57_82));
	PE pe57_83(.x(x83),.w(w57_82),.acc(r57_82),.res(r57_83),.clk(clk),.wout(w57_83));
	PE pe57_84(.x(x84),.w(w57_83),.acc(r57_83),.res(r57_84),.clk(clk),.wout(w57_84));
	PE pe57_85(.x(x85),.w(w57_84),.acc(r57_84),.res(r57_85),.clk(clk),.wout(w57_85));
	PE pe57_86(.x(x86),.w(w57_85),.acc(r57_85),.res(r57_86),.clk(clk),.wout(w57_86));
	PE pe57_87(.x(x87),.w(w57_86),.acc(r57_86),.res(r57_87),.clk(clk),.wout(w57_87));
	PE pe57_88(.x(x88),.w(w57_87),.acc(r57_87),.res(r57_88),.clk(clk),.wout(w57_88));
	PE pe57_89(.x(x89),.w(w57_88),.acc(r57_88),.res(r57_89),.clk(clk),.wout(w57_89));
	PE pe57_90(.x(x90),.w(w57_89),.acc(r57_89),.res(r57_90),.clk(clk),.wout(w57_90));
	PE pe57_91(.x(x91),.w(w57_90),.acc(r57_90),.res(r57_91),.clk(clk),.wout(w57_91));
	PE pe57_92(.x(x92),.w(w57_91),.acc(r57_91),.res(r57_92),.clk(clk),.wout(w57_92));
	PE pe57_93(.x(x93),.w(w57_92),.acc(r57_92),.res(r57_93),.clk(clk),.wout(w57_93));
	PE pe57_94(.x(x94),.w(w57_93),.acc(r57_93),.res(r57_94),.clk(clk),.wout(w57_94));
	PE pe57_95(.x(x95),.w(w57_94),.acc(r57_94),.res(r57_95),.clk(clk),.wout(w57_95));
	PE pe57_96(.x(x96),.w(w57_95),.acc(r57_95),.res(r57_96),.clk(clk),.wout(w57_96));
	PE pe57_97(.x(x97),.w(w57_96),.acc(r57_96),.res(r57_97),.clk(clk),.wout(w57_97));
	PE pe57_98(.x(x98),.w(w57_97),.acc(r57_97),.res(r57_98),.clk(clk),.wout(w57_98));
	PE pe57_99(.x(x99),.w(w57_98),.acc(r57_98),.res(r57_99),.clk(clk),.wout(w57_99));
	PE pe57_100(.x(x100),.w(w57_99),.acc(r57_99),.res(r57_100),.clk(clk),.wout(w57_100));
	PE pe57_101(.x(x101),.w(w57_100),.acc(r57_100),.res(r57_101),.clk(clk),.wout(w57_101));
	PE pe57_102(.x(x102),.w(w57_101),.acc(r57_101),.res(r57_102),.clk(clk),.wout(w57_102));
	PE pe57_103(.x(x103),.w(w57_102),.acc(r57_102),.res(r57_103),.clk(clk),.wout(w57_103));
	PE pe57_104(.x(x104),.w(w57_103),.acc(r57_103),.res(r57_104),.clk(clk),.wout(w57_104));
	PE pe57_105(.x(x105),.w(w57_104),.acc(r57_104),.res(r57_105),.clk(clk),.wout(w57_105));
	PE pe57_106(.x(x106),.w(w57_105),.acc(r57_105),.res(r57_106),.clk(clk),.wout(w57_106));
	PE pe57_107(.x(x107),.w(w57_106),.acc(r57_106),.res(r57_107),.clk(clk),.wout(w57_107));
	PE pe57_108(.x(x108),.w(w57_107),.acc(r57_107),.res(r57_108),.clk(clk),.wout(w57_108));
	PE pe57_109(.x(x109),.w(w57_108),.acc(r57_108),.res(r57_109),.clk(clk),.wout(w57_109));
	PE pe57_110(.x(x110),.w(w57_109),.acc(r57_109),.res(r57_110),.clk(clk),.wout(w57_110));
	PE pe57_111(.x(x111),.w(w57_110),.acc(r57_110),.res(r57_111),.clk(clk),.wout(w57_111));
	PE pe57_112(.x(x112),.w(w57_111),.acc(r57_111),.res(r57_112),.clk(clk),.wout(w57_112));
	PE pe57_113(.x(x113),.w(w57_112),.acc(r57_112),.res(r57_113),.clk(clk),.wout(w57_113));
	PE pe57_114(.x(x114),.w(w57_113),.acc(r57_113),.res(r57_114),.clk(clk),.wout(w57_114));
	PE pe57_115(.x(x115),.w(w57_114),.acc(r57_114),.res(r57_115),.clk(clk),.wout(w57_115));
	PE pe57_116(.x(x116),.w(w57_115),.acc(r57_115),.res(r57_116),.clk(clk),.wout(w57_116));
	PE pe57_117(.x(x117),.w(w57_116),.acc(r57_116),.res(r57_117),.clk(clk),.wout(w57_117));
	PE pe57_118(.x(x118),.w(w57_117),.acc(r57_117),.res(r57_118),.clk(clk),.wout(w57_118));
	PE pe57_119(.x(x119),.w(w57_118),.acc(r57_118),.res(r57_119),.clk(clk),.wout(w57_119));
	PE pe57_120(.x(x120),.w(w57_119),.acc(r57_119),.res(r57_120),.clk(clk),.wout(w57_120));
	PE pe57_121(.x(x121),.w(w57_120),.acc(r57_120),.res(r57_121),.clk(clk),.wout(w57_121));
	PE pe57_122(.x(x122),.w(w57_121),.acc(r57_121),.res(r57_122),.clk(clk),.wout(w57_122));
	PE pe57_123(.x(x123),.w(w57_122),.acc(r57_122),.res(r57_123),.clk(clk),.wout(w57_123));
	PE pe57_124(.x(x124),.w(w57_123),.acc(r57_123),.res(r57_124),.clk(clk),.wout(w57_124));
	PE pe57_125(.x(x125),.w(w57_124),.acc(r57_124),.res(r57_125),.clk(clk),.wout(w57_125));
	PE pe57_126(.x(x126),.w(w57_125),.acc(r57_125),.res(r57_126),.clk(clk),.wout(w57_126));
	PE pe57_127(.x(x127),.w(w57_126),.acc(r57_126),.res(result57),.clk(clk),.wout(weight57));

	PE pe58_0(.x(x0),.w(w58),.acc(32'h0),.res(r58_0),.clk(clk),.wout(w58_0));
	PE pe58_1(.x(x1),.w(w58_0),.acc(r58_0),.res(r58_1),.clk(clk),.wout(w58_1));
	PE pe58_2(.x(x2),.w(w58_1),.acc(r58_1),.res(r58_2),.clk(clk),.wout(w58_2));
	PE pe58_3(.x(x3),.w(w58_2),.acc(r58_2),.res(r58_3),.clk(clk),.wout(w58_3));
	PE pe58_4(.x(x4),.w(w58_3),.acc(r58_3),.res(r58_4),.clk(clk),.wout(w58_4));
	PE pe58_5(.x(x5),.w(w58_4),.acc(r58_4),.res(r58_5),.clk(clk),.wout(w58_5));
	PE pe58_6(.x(x6),.w(w58_5),.acc(r58_5),.res(r58_6),.clk(clk),.wout(w58_6));
	PE pe58_7(.x(x7),.w(w58_6),.acc(r58_6),.res(r58_7),.clk(clk),.wout(w58_7));
	PE pe58_8(.x(x8),.w(w58_7),.acc(r58_7),.res(r58_8),.clk(clk),.wout(w58_8));
	PE pe58_9(.x(x9),.w(w58_8),.acc(r58_8),.res(r58_9),.clk(clk),.wout(w58_9));
	PE pe58_10(.x(x10),.w(w58_9),.acc(r58_9),.res(r58_10),.clk(clk),.wout(w58_10));
	PE pe58_11(.x(x11),.w(w58_10),.acc(r58_10),.res(r58_11),.clk(clk),.wout(w58_11));
	PE pe58_12(.x(x12),.w(w58_11),.acc(r58_11),.res(r58_12),.clk(clk),.wout(w58_12));
	PE pe58_13(.x(x13),.w(w58_12),.acc(r58_12),.res(r58_13),.clk(clk),.wout(w58_13));
	PE pe58_14(.x(x14),.w(w58_13),.acc(r58_13),.res(r58_14),.clk(clk),.wout(w58_14));
	PE pe58_15(.x(x15),.w(w58_14),.acc(r58_14),.res(r58_15),.clk(clk),.wout(w58_15));
	PE pe58_16(.x(x16),.w(w58_15),.acc(r58_15),.res(r58_16),.clk(clk),.wout(w58_16));
	PE pe58_17(.x(x17),.w(w58_16),.acc(r58_16),.res(r58_17),.clk(clk),.wout(w58_17));
	PE pe58_18(.x(x18),.w(w58_17),.acc(r58_17),.res(r58_18),.clk(clk),.wout(w58_18));
	PE pe58_19(.x(x19),.w(w58_18),.acc(r58_18),.res(r58_19),.clk(clk),.wout(w58_19));
	PE pe58_20(.x(x20),.w(w58_19),.acc(r58_19),.res(r58_20),.clk(clk),.wout(w58_20));
	PE pe58_21(.x(x21),.w(w58_20),.acc(r58_20),.res(r58_21),.clk(clk),.wout(w58_21));
	PE pe58_22(.x(x22),.w(w58_21),.acc(r58_21),.res(r58_22),.clk(clk),.wout(w58_22));
	PE pe58_23(.x(x23),.w(w58_22),.acc(r58_22),.res(r58_23),.clk(clk),.wout(w58_23));
	PE pe58_24(.x(x24),.w(w58_23),.acc(r58_23),.res(r58_24),.clk(clk),.wout(w58_24));
	PE pe58_25(.x(x25),.w(w58_24),.acc(r58_24),.res(r58_25),.clk(clk),.wout(w58_25));
	PE pe58_26(.x(x26),.w(w58_25),.acc(r58_25),.res(r58_26),.clk(clk),.wout(w58_26));
	PE pe58_27(.x(x27),.w(w58_26),.acc(r58_26),.res(r58_27),.clk(clk),.wout(w58_27));
	PE pe58_28(.x(x28),.w(w58_27),.acc(r58_27),.res(r58_28),.clk(clk),.wout(w58_28));
	PE pe58_29(.x(x29),.w(w58_28),.acc(r58_28),.res(r58_29),.clk(clk),.wout(w58_29));
	PE pe58_30(.x(x30),.w(w58_29),.acc(r58_29),.res(r58_30),.clk(clk),.wout(w58_30));
	PE pe58_31(.x(x31),.w(w58_30),.acc(r58_30),.res(r58_31),.clk(clk),.wout(w58_31));
	PE pe58_32(.x(x32),.w(w58_31),.acc(r58_31),.res(r58_32),.clk(clk),.wout(w58_32));
	PE pe58_33(.x(x33),.w(w58_32),.acc(r58_32),.res(r58_33),.clk(clk),.wout(w58_33));
	PE pe58_34(.x(x34),.w(w58_33),.acc(r58_33),.res(r58_34),.clk(clk),.wout(w58_34));
	PE pe58_35(.x(x35),.w(w58_34),.acc(r58_34),.res(r58_35),.clk(clk),.wout(w58_35));
	PE pe58_36(.x(x36),.w(w58_35),.acc(r58_35),.res(r58_36),.clk(clk),.wout(w58_36));
	PE pe58_37(.x(x37),.w(w58_36),.acc(r58_36),.res(r58_37),.clk(clk),.wout(w58_37));
	PE pe58_38(.x(x38),.w(w58_37),.acc(r58_37),.res(r58_38),.clk(clk),.wout(w58_38));
	PE pe58_39(.x(x39),.w(w58_38),.acc(r58_38),.res(r58_39),.clk(clk),.wout(w58_39));
	PE pe58_40(.x(x40),.w(w58_39),.acc(r58_39),.res(r58_40),.clk(clk),.wout(w58_40));
	PE pe58_41(.x(x41),.w(w58_40),.acc(r58_40),.res(r58_41),.clk(clk),.wout(w58_41));
	PE pe58_42(.x(x42),.w(w58_41),.acc(r58_41),.res(r58_42),.clk(clk),.wout(w58_42));
	PE pe58_43(.x(x43),.w(w58_42),.acc(r58_42),.res(r58_43),.clk(clk),.wout(w58_43));
	PE pe58_44(.x(x44),.w(w58_43),.acc(r58_43),.res(r58_44),.clk(clk),.wout(w58_44));
	PE pe58_45(.x(x45),.w(w58_44),.acc(r58_44),.res(r58_45),.clk(clk),.wout(w58_45));
	PE pe58_46(.x(x46),.w(w58_45),.acc(r58_45),.res(r58_46),.clk(clk),.wout(w58_46));
	PE pe58_47(.x(x47),.w(w58_46),.acc(r58_46),.res(r58_47),.clk(clk),.wout(w58_47));
	PE pe58_48(.x(x48),.w(w58_47),.acc(r58_47),.res(r58_48),.clk(clk),.wout(w58_48));
	PE pe58_49(.x(x49),.w(w58_48),.acc(r58_48),.res(r58_49),.clk(clk),.wout(w58_49));
	PE pe58_50(.x(x50),.w(w58_49),.acc(r58_49),.res(r58_50),.clk(clk),.wout(w58_50));
	PE pe58_51(.x(x51),.w(w58_50),.acc(r58_50),.res(r58_51),.clk(clk),.wout(w58_51));
	PE pe58_52(.x(x52),.w(w58_51),.acc(r58_51),.res(r58_52),.clk(clk),.wout(w58_52));
	PE pe58_53(.x(x53),.w(w58_52),.acc(r58_52),.res(r58_53),.clk(clk),.wout(w58_53));
	PE pe58_54(.x(x54),.w(w58_53),.acc(r58_53),.res(r58_54),.clk(clk),.wout(w58_54));
	PE pe58_55(.x(x55),.w(w58_54),.acc(r58_54),.res(r58_55),.clk(clk),.wout(w58_55));
	PE pe58_56(.x(x56),.w(w58_55),.acc(r58_55),.res(r58_56),.clk(clk),.wout(w58_56));
	PE pe58_57(.x(x57),.w(w58_56),.acc(r58_56),.res(r58_57),.clk(clk),.wout(w58_57));
	PE pe58_58(.x(x58),.w(w58_57),.acc(r58_57),.res(r58_58),.clk(clk),.wout(w58_58));
	PE pe58_59(.x(x59),.w(w58_58),.acc(r58_58),.res(r58_59),.clk(clk),.wout(w58_59));
	PE pe58_60(.x(x60),.w(w58_59),.acc(r58_59),.res(r58_60),.clk(clk),.wout(w58_60));
	PE pe58_61(.x(x61),.w(w58_60),.acc(r58_60),.res(r58_61),.clk(clk),.wout(w58_61));
	PE pe58_62(.x(x62),.w(w58_61),.acc(r58_61),.res(r58_62),.clk(clk),.wout(w58_62));
	PE pe58_63(.x(x63),.w(w58_62),.acc(r58_62),.res(r58_63),.clk(clk),.wout(w58_63));
	PE pe58_64(.x(x64),.w(w58_63),.acc(r58_63),.res(r58_64),.clk(clk),.wout(w58_64));
	PE pe58_65(.x(x65),.w(w58_64),.acc(r58_64),.res(r58_65),.clk(clk),.wout(w58_65));
	PE pe58_66(.x(x66),.w(w58_65),.acc(r58_65),.res(r58_66),.clk(clk),.wout(w58_66));
	PE pe58_67(.x(x67),.w(w58_66),.acc(r58_66),.res(r58_67),.clk(clk),.wout(w58_67));
	PE pe58_68(.x(x68),.w(w58_67),.acc(r58_67),.res(r58_68),.clk(clk),.wout(w58_68));
	PE pe58_69(.x(x69),.w(w58_68),.acc(r58_68),.res(r58_69),.clk(clk),.wout(w58_69));
	PE pe58_70(.x(x70),.w(w58_69),.acc(r58_69),.res(r58_70),.clk(clk),.wout(w58_70));
	PE pe58_71(.x(x71),.w(w58_70),.acc(r58_70),.res(r58_71),.clk(clk),.wout(w58_71));
	PE pe58_72(.x(x72),.w(w58_71),.acc(r58_71),.res(r58_72),.clk(clk),.wout(w58_72));
	PE pe58_73(.x(x73),.w(w58_72),.acc(r58_72),.res(r58_73),.clk(clk),.wout(w58_73));
	PE pe58_74(.x(x74),.w(w58_73),.acc(r58_73),.res(r58_74),.clk(clk),.wout(w58_74));
	PE pe58_75(.x(x75),.w(w58_74),.acc(r58_74),.res(r58_75),.clk(clk),.wout(w58_75));
	PE pe58_76(.x(x76),.w(w58_75),.acc(r58_75),.res(r58_76),.clk(clk),.wout(w58_76));
	PE pe58_77(.x(x77),.w(w58_76),.acc(r58_76),.res(r58_77),.clk(clk),.wout(w58_77));
	PE pe58_78(.x(x78),.w(w58_77),.acc(r58_77),.res(r58_78),.clk(clk),.wout(w58_78));
	PE pe58_79(.x(x79),.w(w58_78),.acc(r58_78),.res(r58_79),.clk(clk),.wout(w58_79));
	PE pe58_80(.x(x80),.w(w58_79),.acc(r58_79),.res(r58_80),.clk(clk),.wout(w58_80));
	PE pe58_81(.x(x81),.w(w58_80),.acc(r58_80),.res(r58_81),.clk(clk),.wout(w58_81));
	PE pe58_82(.x(x82),.w(w58_81),.acc(r58_81),.res(r58_82),.clk(clk),.wout(w58_82));
	PE pe58_83(.x(x83),.w(w58_82),.acc(r58_82),.res(r58_83),.clk(clk),.wout(w58_83));
	PE pe58_84(.x(x84),.w(w58_83),.acc(r58_83),.res(r58_84),.clk(clk),.wout(w58_84));
	PE pe58_85(.x(x85),.w(w58_84),.acc(r58_84),.res(r58_85),.clk(clk),.wout(w58_85));
	PE pe58_86(.x(x86),.w(w58_85),.acc(r58_85),.res(r58_86),.clk(clk),.wout(w58_86));
	PE pe58_87(.x(x87),.w(w58_86),.acc(r58_86),.res(r58_87),.clk(clk),.wout(w58_87));
	PE pe58_88(.x(x88),.w(w58_87),.acc(r58_87),.res(r58_88),.clk(clk),.wout(w58_88));
	PE pe58_89(.x(x89),.w(w58_88),.acc(r58_88),.res(r58_89),.clk(clk),.wout(w58_89));
	PE pe58_90(.x(x90),.w(w58_89),.acc(r58_89),.res(r58_90),.clk(clk),.wout(w58_90));
	PE pe58_91(.x(x91),.w(w58_90),.acc(r58_90),.res(r58_91),.clk(clk),.wout(w58_91));
	PE pe58_92(.x(x92),.w(w58_91),.acc(r58_91),.res(r58_92),.clk(clk),.wout(w58_92));
	PE pe58_93(.x(x93),.w(w58_92),.acc(r58_92),.res(r58_93),.clk(clk),.wout(w58_93));
	PE pe58_94(.x(x94),.w(w58_93),.acc(r58_93),.res(r58_94),.clk(clk),.wout(w58_94));
	PE pe58_95(.x(x95),.w(w58_94),.acc(r58_94),.res(r58_95),.clk(clk),.wout(w58_95));
	PE pe58_96(.x(x96),.w(w58_95),.acc(r58_95),.res(r58_96),.clk(clk),.wout(w58_96));
	PE pe58_97(.x(x97),.w(w58_96),.acc(r58_96),.res(r58_97),.clk(clk),.wout(w58_97));
	PE pe58_98(.x(x98),.w(w58_97),.acc(r58_97),.res(r58_98),.clk(clk),.wout(w58_98));
	PE pe58_99(.x(x99),.w(w58_98),.acc(r58_98),.res(r58_99),.clk(clk),.wout(w58_99));
	PE pe58_100(.x(x100),.w(w58_99),.acc(r58_99),.res(r58_100),.clk(clk),.wout(w58_100));
	PE pe58_101(.x(x101),.w(w58_100),.acc(r58_100),.res(r58_101),.clk(clk),.wout(w58_101));
	PE pe58_102(.x(x102),.w(w58_101),.acc(r58_101),.res(r58_102),.clk(clk),.wout(w58_102));
	PE pe58_103(.x(x103),.w(w58_102),.acc(r58_102),.res(r58_103),.clk(clk),.wout(w58_103));
	PE pe58_104(.x(x104),.w(w58_103),.acc(r58_103),.res(r58_104),.clk(clk),.wout(w58_104));
	PE pe58_105(.x(x105),.w(w58_104),.acc(r58_104),.res(r58_105),.clk(clk),.wout(w58_105));
	PE pe58_106(.x(x106),.w(w58_105),.acc(r58_105),.res(r58_106),.clk(clk),.wout(w58_106));
	PE pe58_107(.x(x107),.w(w58_106),.acc(r58_106),.res(r58_107),.clk(clk),.wout(w58_107));
	PE pe58_108(.x(x108),.w(w58_107),.acc(r58_107),.res(r58_108),.clk(clk),.wout(w58_108));
	PE pe58_109(.x(x109),.w(w58_108),.acc(r58_108),.res(r58_109),.clk(clk),.wout(w58_109));
	PE pe58_110(.x(x110),.w(w58_109),.acc(r58_109),.res(r58_110),.clk(clk),.wout(w58_110));
	PE pe58_111(.x(x111),.w(w58_110),.acc(r58_110),.res(r58_111),.clk(clk),.wout(w58_111));
	PE pe58_112(.x(x112),.w(w58_111),.acc(r58_111),.res(r58_112),.clk(clk),.wout(w58_112));
	PE pe58_113(.x(x113),.w(w58_112),.acc(r58_112),.res(r58_113),.clk(clk),.wout(w58_113));
	PE pe58_114(.x(x114),.w(w58_113),.acc(r58_113),.res(r58_114),.clk(clk),.wout(w58_114));
	PE pe58_115(.x(x115),.w(w58_114),.acc(r58_114),.res(r58_115),.clk(clk),.wout(w58_115));
	PE pe58_116(.x(x116),.w(w58_115),.acc(r58_115),.res(r58_116),.clk(clk),.wout(w58_116));
	PE pe58_117(.x(x117),.w(w58_116),.acc(r58_116),.res(r58_117),.clk(clk),.wout(w58_117));
	PE pe58_118(.x(x118),.w(w58_117),.acc(r58_117),.res(r58_118),.clk(clk),.wout(w58_118));
	PE pe58_119(.x(x119),.w(w58_118),.acc(r58_118),.res(r58_119),.clk(clk),.wout(w58_119));
	PE pe58_120(.x(x120),.w(w58_119),.acc(r58_119),.res(r58_120),.clk(clk),.wout(w58_120));
	PE pe58_121(.x(x121),.w(w58_120),.acc(r58_120),.res(r58_121),.clk(clk),.wout(w58_121));
	PE pe58_122(.x(x122),.w(w58_121),.acc(r58_121),.res(r58_122),.clk(clk),.wout(w58_122));
	PE pe58_123(.x(x123),.w(w58_122),.acc(r58_122),.res(r58_123),.clk(clk),.wout(w58_123));
	PE pe58_124(.x(x124),.w(w58_123),.acc(r58_123),.res(r58_124),.clk(clk),.wout(w58_124));
	PE pe58_125(.x(x125),.w(w58_124),.acc(r58_124),.res(r58_125),.clk(clk),.wout(w58_125));
	PE pe58_126(.x(x126),.w(w58_125),.acc(r58_125),.res(r58_126),.clk(clk),.wout(w58_126));
	PE pe58_127(.x(x127),.w(w58_126),.acc(r58_126),.res(result58),.clk(clk),.wout(weight58));

	PE pe59_0(.x(x0),.w(w59),.acc(32'h0),.res(r59_0),.clk(clk),.wout(w59_0));
	PE pe59_1(.x(x1),.w(w59_0),.acc(r59_0),.res(r59_1),.clk(clk),.wout(w59_1));
	PE pe59_2(.x(x2),.w(w59_1),.acc(r59_1),.res(r59_2),.clk(clk),.wout(w59_2));
	PE pe59_3(.x(x3),.w(w59_2),.acc(r59_2),.res(r59_3),.clk(clk),.wout(w59_3));
	PE pe59_4(.x(x4),.w(w59_3),.acc(r59_3),.res(r59_4),.clk(clk),.wout(w59_4));
	PE pe59_5(.x(x5),.w(w59_4),.acc(r59_4),.res(r59_5),.clk(clk),.wout(w59_5));
	PE pe59_6(.x(x6),.w(w59_5),.acc(r59_5),.res(r59_6),.clk(clk),.wout(w59_6));
	PE pe59_7(.x(x7),.w(w59_6),.acc(r59_6),.res(r59_7),.clk(clk),.wout(w59_7));
	PE pe59_8(.x(x8),.w(w59_7),.acc(r59_7),.res(r59_8),.clk(clk),.wout(w59_8));
	PE pe59_9(.x(x9),.w(w59_8),.acc(r59_8),.res(r59_9),.clk(clk),.wout(w59_9));
	PE pe59_10(.x(x10),.w(w59_9),.acc(r59_9),.res(r59_10),.clk(clk),.wout(w59_10));
	PE pe59_11(.x(x11),.w(w59_10),.acc(r59_10),.res(r59_11),.clk(clk),.wout(w59_11));
	PE pe59_12(.x(x12),.w(w59_11),.acc(r59_11),.res(r59_12),.clk(clk),.wout(w59_12));
	PE pe59_13(.x(x13),.w(w59_12),.acc(r59_12),.res(r59_13),.clk(clk),.wout(w59_13));
	PE pe59_14(.x(x14),.w(w59_13),.acc(r59_13),.res(r59_14),.clk(clk),.wout(w59_14));
	PE pe59_15(.x(x15),.w(w59_14),.acc(r59_14),.res(r59_15),.clk(clk),.wout(w59_15));
	PE pe59_16(.x(x16),.w(w59_15),.acc(r59_15),.res(r59_16),.clk(clk),.wout(w59_16));
	PE pe59_17(.x(x17),.w(w59_16),.acc(r59_16),.res(r59_17),.clk(clk),.wout(w59_17));
	PE pe59_18(.x(x18),.w(w59_17),.acc(r59_17),.res(r59_18),.clk(clk),.wout(w59_18));
	PE pe59_19(.x(x19),.w(w59_18),.acc(r59_18),.res(r59_19),.clk(clk),.wout(w59_19));
	PE pe59_20(.x(x20),.w(w59_19),.acc(r59_19),.res(r59_20),.clk(clk),.wout(w59_20));
	PE pe59_21(.x(x21),.w(w59_20),.acc(r59_20),.res(r59_21),.clk(clk),.wout(w59_21));
	PE pe59_22(.x(x22),.w(w59_21),.acc(r59_21),.res(r59_22),.clk(clk),.wout(w59_22));
	PE pe59_23(.x(x23),.w(w59_22),.acc(r59_22),.res(r59_23),.clk(clk),.wout(w59_23));
	PE pe59_24(.x(x24),.w(w59_23),.acc(r59_23),.res(r59_24),.clk(clk),.wout(w59_24));
	PE pe59_25(.x(x25),.w(w59_24),.acc(r59_24),.res(r59_25),.clk(clk),.wout(w59_25));
	PE pe59_26(.x(x26),.w(w59_25),.acc(r59_25),.res(r59_26),.clk(clk),.wout(w59_26));
	PE pe59_27(.x(x27),.w(w59_26),.acc(r59_26),.res(r59_27),.clk(clk),.wout(w59_27));
	PE pe59_28(.x(x28),.w(w59_27),.acc(r59_27),.res(r59_28),.clk(clk),.wout(w59_28));
	PE pe59_29(.x(x29),.w(w59_28),.acc(r59_28),.res(r59_29),.clk(clk),.wout(w59_29));
	PE pe59_30(.x(x30),.w(w59_29),.acc(r59_29),.res(r59_30),.clk(clk),.wout(w59_30));
	PE pe59_31(.x(x31),.w(w59_30),.acc(r59_30),.res(r59_31),.clk(clk),.wout(w59_31));
	PE pe59_32(.x(x32),.w(w59_31),.acc(r59_31),.res(r59_32),.clk(clk),.wout(w59_32));
	PE pe59_33(.x(x33),.w(w59_32),.acc(r59_32),.res(r59_33),.clk(clk),.wout(w59_33));
	PE pe59_34(.x(x34),.w(w59_33),.acc(r59_33),.res(r59_34),.clk(clk),.wout(w59_34));
	PE pe59_35(.x(x35),.w(w59_34),.acc(r59_34),.res(r59_35),.clk(clk),.wout(w59_35));
	PE pe59_36(.x(x36),.w(w59_35),.acc(r59_35),.res(r59_36),.clk(clk),.wout(w59_36));
	PE pe59_37(.x(x37),.w(w59_36),.acc(r59_36),.res(r59_37),.clk(clk),.wout(w59_37));
	PE pe59_38(.x(x38),.w(w59_37),.acc(r59_37),.res(r59_38),.clk(clk),.wout(w59_38));
	PE pe59_39(.x(x39),.w(w59_38),.acc(r59_38),.res(r59_39),.clk(clk),.wout(w59_39));
	PE pe59_40(.x(x40),.w(w59_39),.acc(r59_39),.res(r59_40),.clk(clk),.wout(w59_40));
	PE pe59_41(.x(x41),.w(w59_40),.acc(r59_40),.res(r59_41),.clk(clk),.wout(w59_41));
	PE pe59_42(.x(x42),.w(w59_41),.acc(r59_41),.res(r59_42),.clk(clk),.wout(w59_42));
	PE pe59_43(.x(x43),.w(w59_42),.acc(r59_42),.res(r59_43),.clk(clk),.wout(w59_43));
	PE pe59_44(.x(x44),.w(w59_43),.acc(r59_43),.res(r59_44),.clk(clk),.wout(w59_44));
	PE pe59_45(.x(x45),.w(w59_44),.acc(r59_44),.res(r59_45),.clk(clk),.wout(w59_45));
	PE pe59_46(.x(x46),.w(w59_45),.acc(r59_45),.res(r59_46),.clk(clk),.wout(w59_46));
	PE pe59_47(.x(x47),.w(w59_46),.acc(r59_46),.res(r59_47),.clk(clk),.wout(w59_47));
	PE pe59_48(.x(x48),.w(w59_47),.acc(r59_47),.res(r59_48),.clk(clk),.wout(w59_48));
	PE pe59_49(.x(x49),.w(w59_48),.acc(r59_48),.res(r59_49),.clk(clk),.wout(w59_49));
	PE pe59_50(.x(x50),.w(w59_49),.acc(r59_49),.res(r59_50),.clk(clk),.wout(w59_50));
	PE pe59_51(.x(x51),.w(w59_50),.acc(r59_50),.res(r59_51),.clk(clk),.wout(w59_51));
	PE pe59_52(.x(x52),.w(w59_51),.acc(r59_51),.res(r59_52),.clk(clk),.wout(w59_52));
	PE pe59_53(.x(x53),.w(w59_52),.acc(r59_52),.res(r59_53),.clk(clk),.wout(w59_53));
	PE pe59_54(.x(x54),.w(w59_53),.acc(r59_53),.res(r59_54),.clk(clk),.wout(w59_54));
	PE pe59_55(.x(x55),.w(w59_54),.acc(r59_54),.res(r59_55),.clk(clk),.wout(w59_55));
	PE pe59_56(.x(x56),.w(w59_55),.acc(r59_55),.res(r59_56),.clk(clk),.wout(w59_56));
	PE pe59_57(.x(x57),.w(w59_56),.acc(r59_56),.res(r59_57),.clk(clk),.wout(w59_57));
	PE pe59_58(.x(x58),.w(w59_57),.acc(r59_57),.res(r59_58),.clk(clk),.wout(w59_58));
	PE pe59_59(.x(x59),.w(w59_58),.acc(r59_58),.res(r59_59),.clk(clk),.wout(w59_59));
	PE pe59_60(.x(x60),.w(w59_59),.acc(r59_59),.res(r59_60),.clk(clk),.wout(w59_60));
	PE pe59_61(.x(x61),.w(w59_60),.acc(r59_60),.res(r59_61),.clk(clk),.wout(w59_61));
	PE pe59_62(.x(x62),.w(w59_61),.acc(r59_61),.res(r59_62),.clk(clk),.wout(w59_62));
	PE pe59_63(.x(x63),.w(w59_62),.acc(r59_62),.res(r59_63),.clk(clk),.wout(w59_63));
	PE pe59_64(.x(x64),.w(w59_63),.acc(r59_63),.res(r59_64),.clk(clk),.wout(w59_64));
	PE pe59_65(.x(x65),.w(w59_64),.acc(r59_64),.res(r59_65),.clk(clk),.wout(w59_65));
	PE pe59_66(.x(x66),.w(w59_65),.acc(r59_65),.res(r59_66),.clk(clk),.wout(w59_66));
	PE pe59_67(.x(x67),.w(w59_66),.acc(r59_66),.res(r59_67),.clk(clk),.wout(w59_67));
	PE pe59_68(.x(x68),.w(w59_67),.acc(r59_67),.res(r59_68),.clk(clk),.wout(w59_68));
	PE pe59_69(.x(x69),.w(w59_68),.acc(r59_68),.res(r59_69),.clk(clk),.wout(w59_69));
	PE pe59_70(.x(x70),.w(w59_69),.acc(r59_69),.res(r59_70),.clk(clk),.wout(w59_70));
	PE pe59_71(.x(x71),.w(w59_70),.acc(r59_70),.res(r59_71),.clk(clk),.wout(w59_71));
	PE pe59_72(.x(x72),.w(w59_71),.acc(r59_71),.res(r59_72),.clk(clk),.wout(w59_72));
	PE pe59_73(.x(x73),.w(w59_72),.acc(r59_72),.res(r59_73),.clk(clk),.wout(w59_73));
	PE pe59_74(.x(x74),.w(w59_73),.acc(r59_73),.res(r59_74),.clk(clk),.wout(w59_74));
	PE pe59_75(.x(x75),.w(w59_74),.acc(r59_74),.res(r59_75),.clk(clk),.wout(w59_75));
	PE pe59_76(.x(x76),.w(w59_75),.acc(r59_75),.res(r59_76),.clk(clk),.wout(w59_76));
	PE pe59_77(.x(x77),.w(w59_76),.acc(r59_76),.res(r59_77),.clk(clk),.wout(w59_77));
	PE pe59_78(.x(x78),.w(w59_77),.acc(r59_77),.res(r59_78),.clk(clk),.wout(w59_78));
	PE pe59_79(.x(x79),.w(w59_78),.acc(r59_78),.res(r59_79),.clk(clk),.wout(w59_79));
	PE pe59_80(.x(x80),.w(w59_79),.acc(r59_79),.res(r59_80),.clk(clk),.wout(w59_80));
	PE pe59_81(.x(x81),.w(w59_80),.acc(r59_80),.res(r59_81),.clk(clk),.wout(w59_81));
	PE pe59_82(.x(x82),.w(w59_81),.acc(r59_81),.res(r59_82),.clk(clk),.wout(w59_82));
	PE pe59_83(.x(x83),.w(w59_82),.acc(r59_82),.res(r59_83),.clk(clk),.wout(w59_83));
	PE pe59_84(.x(x84),.w(w59_83),.acc(r59_83),.res(r59_84),.clk(clk),.wout(w59_84));
	PE pe59_85(.x(x85),.w(w59_84),.acc(r59_84),.res(r59_85),.clk(clk),.wout(w59_85));
	PE pe59_86(.x(x86),.w(w59_85),.acc(r59_85),.res(r59_86),.clk(clk),.wout(w59_86));
	PE pe59_87(.x(x87),.w(w59_86),.acc(r59_86),.res(r59_87),.clk(clk),.wout(w59_87));
	PE pe59_88(.x(x88),.w(w59_87),.acc(r59_87),.res(r59_88),.clk(clk),.wout(w59_88));
	PE pe59_89(.x(x89),.w(w59_88),.acc(r59_88),.res(r59_89),.clk(clk),.wout(w59_89));
	PE pe59_90(.x(x90),.w(w59_89),.acc(r59_89),.res(r59_90),.clk(clk),.wout(w59_90));
	PE pe59_91(.x(x91),.w(w59_90),.acc(r59_90),.res(r59_91),.clk(clk),.wout(w59_91));
	PE pe59_92(.x(x92),.w(w59_91),.acc(r59_91),.res(r59_92),.clk(clk),.wout(w59_92));
	PE pe59_93(.x(x93),.w(w59_92),.acc(r59_92),.res(r59_93),.clk(clk),.wout(w59_93));
	PE pe59_94(.x(x94),.w(w59_93),.acc(r59_93),.res(r59_94),.clk(clk),.wout(w59_94));
	PE pe59_95(.x(x95),.w(w59_94),.acc(r59_94),.res(r59_95),.clk(clk),.wout(w59_95));
	PE pe59_96(.x(x96),.w(w59_95),.acc(r59_95),.res(r59_96),.clk(clk),.wout(w59_96));
	PE pe59_97(.x(x97),.w(w59_96),.acc(r59_96),.res(r59_97),.clk(clk),.wout(w59_97));
	PE pe59_98(.x(x98),.w(w59_97),.acc(r59_97),.res(r59_98),.clk(clk),.wout(w59_98));
	PE pe59_99(.x(x99),.w(w59_98),.acc(r59_98),.res(r59_99),.clk(clk),.wout(w59_99));
	PE pe59_100(.x(x100),.w(w59_99),.acc(r59_99),.res(r59_100),.clk(clk),.wout(w59_100));
	PE pe59_101(.x(x101),.w(w59_100),.acc(r59_100),.res(r59_101),.clk(clk),.wout(w59_101));
	PE pe59_102(.x(x102),.w(w59_101),.acc(r59_101),.res(r59_102),.clk(clk),.wout(w59_102));
	PE pe59_103(.x(x103),.w(w59_102),.acc(r59_102),.res(r59_103),.clk(clk),.wout(w59_103));
	PE pe59_104(.x(x104),.w(w59_103),.acc(r59_103),.res(r59_104),.clk(clk),.wout(w59_104));
	PE pe59_105(.x(x105),.w(w59_104),.acc(r59_104),.res(r59_105),.clk(clk),.wout(w59_105));
	PE pe59_106(.x(x106),.w(w59_105),.acc(r59_105),.res(r59_106),.clk(clk),.wout(w59_106));
	PE pe59_107(.x(x107),.w(w59_106),.acc(r59_106),.res(r59_107),.clk(clk),.wout(w59_107));
	PE pe59_108(.x(x108),.w(w59_107),.acc(r59_107),.res(r59_108),.clk(clk),.wout(w59_108));
	PE pe59_109(.x(x109),.w(w59_108),.acc(r59_108),.res(r59_109),.clk(clk),.wout(w59_109));
	PE pe59_110(.x(x110),.w(w59_109),.acc(r59_109),.res(r59_110),.clk(clk),.wout(w59_110));
	PE pe59_111(.x(x111),.w(w59_110),.acc(r59_110),.res(r59_111),.clk(clk),.wout(w59_111));
	PE pe59_112(.x(x112),.w(w59_111),.acc(r59_111),.res(r59_112),.clk(clk),.wout(w59_112));
	PE pe59_113(.x(x113),.w(w59_112),.acc(r59_112),.res(r59_113),.clk(clk),.wout(w59_113));
	PE pe59_114(.x(x114),.w(w59_113),.acc(r59_113),.res(r59_114),.clk(clk),.wout(w59_114));
	PE pe59_115(.x(x115),.w(w59_114),.acc(r59_114),.res(r59_115),.clk(clk),.wout(w59_115));
	PE pe59_116(.x(x116),.w(w59_115),.acc(r59_115),.res(r59_116),.clk(clk),.wout(w59_116));
	PE pe59_117(.x(x117),.w(w59_116),.acc(r59_116),.res(r59_117),.clk(clk),.wout(w59_117));
	PE pe59_118(.x(x118),.w(w59_117),.acc(r59_117),.res(r59_118),.clk(clk),.wout(w59_118));
	PE pe59_119(.x(x119),.w(w59_118),.acc(r59_118),.res(r59_119),.clk(clk),.wout(w59_119));
	PE pe59_120(.x(x120),.w(w59_119),.acc(r59_119),.res(r59_120),.clk(clk),.wout(w59_120));
	PE pe59_121(.x(x121),.w(w59_120),.acc(r59_120),.res(r59_121),.clk(clk),.wout(w59_121));
	PE pe59_122(.x(x122),.w(w59_121),.acc(r59_121),.res(r59_122),.clk(clk),.wout(w59_122));
	PE pe59_123(.x(x123),.w(w59_122),.acc(r59_122),.res(r59_123),.clk(clk),.wout(w59_123));
	PE pe59_124(.x(x124),.w(w59_123),.acc(r59_123),.res(r59_124),.clk(clk),.wout(w59_124));
	PE pe59_125(.x(x125),.w(w59_124),.acc(r59_124),.res(r59_125),.clk(clk),.wout(w59_125));
	PE pe59_126(.x(x126),.w(w59_125),.acc(r59_125),.res(r59_126),.clk(clk),.wout(w59_126));
	PE pe59_127(.x(x127),.w(w59_126),.acc(r59_126),.res(result59),.clk(clk),.wout(weight59));

	PE pe60_0(.x(x0),.w(w60),.acc(32'h0),.res(r60_0),.clk(clk),.wout(w60_0));
	PE pe60_1(.x(x1),.w(w60_0),.acc(r60_0),.res(r60_1),.clk(clk),.wout(w60_1));
	PE pe60_2(.x(x2),.w(w60_1),.acc(r60_1),.res(r60_2),.clk(clk),.wout(w60_2));
	PE pe60_3(.x(x3),.w(w60_2),.acc(r60_2),.res(r60_3),.clk(clk),.wout(w60_3));
	PE pe60_4(.x(x4),.w(w60_3),.acc(r60_3),.res(r60_4),.clk(clk),.wout(w60_4));
	PE pe60_5(.x(x5),.w(w60_4),.acc(r60_4),.res(r60_5),.clk(clk),.wout(w60_5));
	PE pe60_6(.x(x6),.w(w60_5),.acc(r60_5),.res(r60_6),.clk(clk),.wout(w60_6));
	PE pe60_7(.x(x7),.w(w60_6),.acc(r60_6),.res(r60_7),.clk(clk),.wout(w60_7));
	PE pe60_8(.x(x8),.w(w60_7),.acc(r60_7),.res(r60_8),.clk(clk),.wout(w60_8));
	PE pe60_9(.x(x9),.w(w60_8),.acc(r60_8),.res(r60_9),.clk(clk),.wout(w60_9));
	PE pe60_10(.x(x10),.w(w60_9),.acc(r60_9),.res(r60_10),.clk(clk),.wout(w60_10));
	PE pe60_11(.x(x11),.w(w60_10),.acc(r60_10),.res(r60_11),.clk(clk),.wout(w60_11));
	PE pe60_12(.x(x12),.w(w60_11),.acc(r60_11),.res(r60_12),.clk(clk),.wout(w60_12));
	PE pe60_13(.x(x13),.w(w60_12),.acc(r60_12),.res(r60_13),.clk(clk),.wout(w60_13));
	PE pe60_14(.x(x14),.w(w60_13),.acc(r60_13),.res(r60_14),.clk(clk),.wout(w60_14));
	PE pe60_15(.x(x15),.w(w60_14),.acc(r60_14),.res(r60_15),.clk(clk),.wout(w60_15));
	PE pe60_16(.x(x16),.w(w60_15),.acc(r60_15),.res(r60_16),.clk(clk),.wout(w60_16));
	PE pe60_17(.x(x17),.w(w60_16),.acc(r60_16),.res(r60_17),.clk(clk),.wout(w60_17));
	PE pe60_18(.x(x18),.w(w60_17),.acc(r60_17),.res(r60_18),.clk(clk),.wout(w60_18));
	PE pe60_19(.x(x19),.w(w60_18),.acc(r60_18),.res(r60_19),.clk(clk),.wout(w60_19));
	PE pe60_20(.x(x20),.w(w60_19),.acc(r60_19),.res(r60_20),.clk(clk),.wout(w60_20));
	PE pe60_21(.x(x21),.w(w60_20),.acc(r60_20),.res(r60_21),.clk(clk),.wout(w60_21));
	PE pe60_22(.x(x22),.w(w60_21),.acc(r60_21),.res(r60_22),.clk(clk),.wout(w60_22));
	PE pe60_23(.x(x23),.w(w60_22),.acc(r60_22),.res(r60_23),.clk(clk),.wout(w60_23));
	PE pe60_24(.x(x24),.w(w60_23),.acc(r60_23),.res(r60_24),.clk(clk),.wout(w60_24));
	PE pe60_25(.x(x25),.w(w60_24),.acc(r60_24),.res(r60_25),.clk(clk),.wout(w60_25));
	PE pe60_26(.x(x26),.w(w60_25),.acc(r60_25),.res(r60_26),.clk(clk),.wout(w60_26));
	PE pe60_27(.x(x27),.w(w60_26),.acc(r60_26),.res(r60_27),.clk(clk),.wout(w60_27));
	PE pe60_28(.x(x28),.w(w60_27),.acc(r60_27),.res(r60_28),.clk(clk),.wout(w60_28));
	PE pe60_29(.x(x29),.w(w60_28),.acc(r60_28),.res(r60_29),.clk(clk),.wout(w60_29));
	PE pe60_30(.x(x30),.w(w60_29),.acc(r60_29),.res(r60_30),.clk(clk),.wout(w60_30));
	PE pe60_31(.x(x31),.w(w60_30),.acc(r60_30),.res(r60_31),.clk(clk),.wout(w60_31));
	PE pe60_32(.x(x32),.w(w60_31),.acc(r60_31),.res(r60_32),.clk(clk),.wout(w60_32));
	PE pe60_33(.x(x33),.w(w60_32),.acc(r60_32),.res(r60_33),.clk(clk),.wout(w60_33));
	PE pe60_34(.x(x34),.w(w60_33),.acc(r60_33),.res(r60_34),.clk(clk),.wout(w60_34));
	PE pe60_35(.x(x35),.w(w60_34),.acc(r60_34),.res(r60_35),.clk(clk),.wout(w60_35));
	PE pe60_36(.x(x36),.w(w60_35),.acc(r60_35),.res(r60_36),.clk(clk),.wout(w60_36));
	PE pe60_37(.x(x37),.w(w60_36),.acc(r60_36),.res(r60_37),.clk(clk),.wout(w60_37));
	PE pe60_38(.x(x38),.w(w60_37),.acc(r60_37),.res(r60_38),.clk(clk),.wout(w60_38));
	PE pe60_39(.x(x39),.w(w60_38),.acc(r60_38),.res(r60_39),.clk(clk),.wout(w60_39));
	PE pe60_40(.x(x40),.w(w60_39),.acc(r60_39),.res(r60_40),.clk(clk),.wout(w60_40));
	PE pe60_41(.x(x41),.w(w60_40),.acc(r60_40),.res(r60_41),.clk(clk),.wout(w60_41));
	PE pe60_42(.x(x42),.w(w60_41),.acc(r60_41),.res(r60_42),.clk(clk),.wout(w60_42));
	PE pe60_43(.x(x43),.w(w60_42),.acc(r60_42),.res(r60_43),.clk(clk),.wout(w60_43));
	PE pe60_44(.x(x44),.w(w60_43),.acc(r60_43),.res(r60_44),.clk(clk),.wout(w60_44));
	PE pe60_45(.x(x45),.w(w60_44),.acc(r60_44),.res(r60_45),.clk(clk),.wout(w60_45));
	PE pe60_46(.x(x46),.w(w60_45),.acc(r60_45),.res(r60_46),.clk(clk),.wout(w60_46));
	PE pe60_47(.x(x47),.w(w60_46),.acc(r60_46),.res(r60_47),.clk(clk),.wout(w60_47));
	PE pe60_48(.x(x48),.w(w60_47),.acc(r60_47),.res(r60_48),.clk(clk),.wout(w60_48));
	PE pe60_49(.x(x49),.w(w60_48),.acc(r60_48),.res(r60_49),.clk(clk),.wout(w60_49));
	PE pe60_50(.x(x50),.w(w60_49),.acc(r60_49),.res(r60_50),.clk(clk),.wout(w60_50));
	PE pe60_51(.x(x51),.w(w60_50),.acc(r60_50),.res(r60_51),.clk(clk),.wout(w60_51));
	PE pe60_52(.x(x52),.w(w60_51),.acc(r60_51),.res(r60_52),.clk(clk),.wout(w60_52));
	PE pe60_53(.x(x53),.w(w60_52),.acc(r60_52),.res(r60_53),.clk(clk),.wout(w60_53));
	PE pe60_54(.x(x54),.w(w60_53),.acc(r60_53),.res(r60_54),.clk(clk),.wout(w60_54));
	PE pe60_55(.x(x55),.w(w60_54),.acc(r60_54),.res(r60_55),.clk(clk),.wout(w60_55));
	PE pe60_56(.x(x56),.w(w60_55),.acc(r60_55),.res(r60_56),.clk(clk),.wout(w60_56));
	PE pe60_57(.x(x57),.w(w60_56),.acc(r60_56),.res(r60_57),.clk(clk),.wout(w60_57));
	PE pe60_58(.x(x58),.w(w60_57),.acc(r60_57),.res(r60_58),.clk(clk),.wout(w60_58));
	PE pe60_59(.x(x59),.w(w60_58),.acc(r60_58),.res(r60_59),.clk(clk),.wout(w60_59));
	PE pe60_60(.x(x60),.w(w60_59),.acc(r60_59),.res(r60_60),.clk(clk),.wout(w60_60));
	PE pe60_61(.x(x61),.w(w60_60),.acc(r60_60),.res(r60_61),.clk(clk),.wout(w60_61));
	PE pe60_62(.x(x62),.w(w60_61),.acc(r60_61),.res(r60_62),.clk(clk),.wout(w60_62));
	PE pe60_63(.x(x63),.w(w60_62),.acc(r60_62),.res(r60_63),.clk(clk),.wout(w60_63));
	PE pe60_64(.x(x64),.w(w60_63),.acc(r60_63),.res(r60_64),.clk(clk),.wout(w60_64));
	PE pe60_65(.x(x65),.w(w60_64),.acc(r60_64),.res(r60_65),.clk(clk),.wout(w60_65));
	PE pe60_66(.x(x66),.w(w60_65),.acc(r60_65),.res(r60_66),.clk(clk),.wout(w60_66));
	PE pe60_67(.x(x67),.w(w60_66),.acc(r60_66),.res(r60_67),.clk(clk),.wout(w60_67));
	PE pe60_68(.x(x68),.w(w60_67),.acc(r60_67),.res(r60_68),.clk(clk),.wout(w60_68));
	PE pe60_69(.x(x69),.w(w60_68),.acc(r60_68),.res(r60_69),.clk(clk),.wout(w60_69));
	PE pe60_70(.x(x70),.w(w60_69),.acc(r60_69),.res(r60_70),.clk(clk),.wout(w60_70));
	PE pe60_71(.x(x71),.w(w60_70),.acc(r60_70),.res(r60_71),.clk(clk),.wout(w60_71));
	PE pe60_72(.x(x72),.w(w60_71),.acc(r60_71),.res(r60_72),.clk(clk),.wout(w60_72));
	PE pe60_73(.x(x73),.w(w60_72),.acc(r60_72),.res(r60_73),.clk(clk),.wout(w60_73));
	PE pe60_74(.x(x74),.w(w60_73),.acc(r60_73),.res(r60_74),.clk(clk),.wout(w60_74));
	PE pe60_75(.x(x75),.w(w60_74),.acc(r60_74),.res(r60_75),.clk(clk),.wout(w60_75));
	PE pe60_76(.x(x76),.w(w60_75),.acc(r60_75),.res(r60_76),.clk(clk),.wout(w60_76));
	PE pe60_77(.x(x77),.w(w60_76),.acc(r60_76),.res(r60_77),.clk(clk),.wout(w60_77));
	PE pe60_78(.x(x78),.w(w60_77),.acc(r60_77),.res(r60_78),.clk(clk),.wout(w60_78));
	PE pe60_79(.x(x79),.w(w60_78),.acc(r60_78),.res(r60_79),.clk(clk),.wout(w60_79));
	PE pe60_80(.x(x80),.w(w60_79),.acc(r60_79),.res(r60_80),.clk(clk),.wout(w60_80));
	PE pe60_81(.x(x81),.w(w60_80),.acc(r60_80),.res(r60_81),.clk(clk),.wout(w60_81));
	PE pe60_82(.x(x82),.w(w60_81),.acc(r60_81),.res(r60_82),.clk(clk),.wout(w60_82));
	PE pe60_83(.x(x83),.w(w60_82),.acc(r60_82),.res(r60_83),.clk(clk),.wout(w60_83));
	PE pe60_84(.x(x84),.w(w60_83),.acc(r60_83),.res(r60_84),.clk(clk),.wout(w60_84));
	PE pe60_85(.x(x85),.w(w60_84),.acc(r60_84),.res(r60_85),.clk(clk),.wout(w60_85));
	PE pe60_86(.x(x86),.w(w60_85),.acc(r60_85),.res(r60_86),.clk(clk),.wout(w60_86));
	PE pe60_87(.x(x87),.w(w60_86),.acc(r60_86),.res(r60_87),.clk(clk),.wout(w60_87));
	PE pe60_88(.x(x88),.w(w60_87),.acc(r60_87),.res(r60_88),.clk(clk),.wout(w60_88));
	PE pe60_89(.x(x89),.w(w60_88),.acc(r60_88),.res(r60_89),.clk(clk),.wout(w60_89));
	PE pe60_90(.x(x90),.w(w60_89),.acc(r60_89),.res(r60_90),.clk(clk),.wout(w60_90));
	PE pe60_91(.x(x91),.w(w60_90),.acc(r60_90),.res(r60_91),.clk(clk),.wout(w60_91));
	PE pe60_92(.x(x92),.w(w60_91),.acc(r60_91),.res(r60_92),.clk(clk),.wout(w60_92));
	PE pe60_93(.x(x93),.w(w60_92),.acc(r60_92),.res(r60_93),.clk(clk),.wout(w60_93));
	PE pe60_94(.x(x94),.w(w60_93),.acc(r60_93),.res(r60_94),.clk(clk),.wout(w60_94));
	PE pe60_95(.x(x95),.w(w60_94),.acc(r60_94),.res(r60_95),.clk(clk),.wout(w60_95));
	PE pe60_96(.x(x96),.w(w60_95),.acc(r60_95),.res(r60_96),.clk(clk),.wout(w60_96));
	PE pe60_97(.x(x97),.w(w60_96),.acc(r60_96),.res(r60_97),.clk(clk),.wout(w60_97));
	PE pe60_98(.x(x98),.w(w60_97),.acc(r60_97),.res(r60_98),.clk(clk),.wout(w60_98));
	PE pe60_99(.x(x99),.w(w60_98),.acc(r60_98),.res(r60_99),.clk(clk),.wout(w60_99));
	PE pe60_100(.x(x100),.w(w60_99),.acc(r60_99),.res(r60_100),.clk(clk),.wout(w60_100));
	PE pe60_101(.x(x101),.w(w60_100),.acc(r60_100),.res(r60_101),.clk(clk),.wout(w60_101));
	PE pe60_102(.x(x102),.w(w60_101),.acc(r60_101),.res(r60_102),.clk(clk),.wout(w60_102));
	PE pe60_103(.x(x103),.w(w60_102),.acc(r60_102),.res(r60_103),.clk(clk),.wout(w60_103));
	PE pe60_104(.x(x104),.w(w60_103),.acc(r60_103),.res(r60_104),.clk(clk),.wout(w60_104));
	PE pe60_105(.x(x105),.w(w60_104),.acc(r60_104),.res(r60_105),.clk(clk),.wout(w60_105));
	PE pe60_106(.x(x106),.w(w60_105),.acc(r60_105),.res(r60_106),.clk(clk),.wout(w60_106));
	PE pe60_107(.x(x107),.w(w60_106),.acc(r60_106),.res(r60_107),.clk(clk),.wout(w60_107));
	PE pe60_108(.x(x108),.w(w60_107),.acc(r60_107),.res(r60_108),.clk(clk),.wout(w60_108));
	PE pe60_109(.x(x109),.w(w60_108),.acc(r60_108),.res(r60_109),.clk(clk),.wout(w60_109));
	PE pe60_110(.x(x110),.w(w60_109),.acc(r60_109),.res(r60_110),.clk(clk),.wout(w60_110));
	PE pe60_111(.x(x111),.w(w60_110),.acc(r60_110),.res(r60_111),.clk(clk),.wout(w60_111));
	PE pe60_112(.x(x112),.w(w60_111),.acc(r60_111),.res(r60_112),.clk(clk),.wout(w60_112));
	PE pe60_113(.x(x113),.w(w60_112),.acc(r60_112),.res(r60_113),.clk(clk),.wout(w60_113));
	PE pe60_114(.x(x114),.w(w60_113),.acc(r60_113),.res(r60_114),.clk(clk),.wout(w60_114));
	PE pe60_115(.x(x115),.w(w60_114),.acc(r60_114),.res(r60_115),.clk(clk),.wout(w60_115));
	PE pe60_116(.x(x116),.w(w60_115),.acc(r60_115),.res(r60_116),.clk(clk),.wout(w60_116));
	PE pe60_117(.x(x117),.w(w60_116),.acc(r60_116),.res(r60_117),.clk(clk),.wout(w60_117));
	PE pe60_118(.x(x118),.w(w60_117),.acc(r60_117),.res(r60_118),.clk(clk),.wout(w60_118));
	PE pe60_119(.x(x119),.w(w60_118),.acc(r60_118),.res(r60_119),.clk(clk),.wout(w60_119));
	PE pe60_120(.x(x120),.w(w60_119),.acc(r60_119),.res(r60_120),.clk(clk),.wout(w60_120));
	PE pe60_121(.x(x121),.w(w60_120),.acc(r60_120),.res(r60_121),.clk(clk),.wout(w60_121));
	PE pe60_122(.x(x122),.w(w60_121),.acc(r60_121),.res(r60_122),.clk(clk),.wout(w60_122));
	PE pe60_123(.x(x123),.w(w60_122),.acc(r60_122),.res(r60_123),.clk(clk),.wout(w60_123));
	PE pe60_124(.x(x124),.w(w60_123),.acc(r60_123),.res(r60_124),.clk(clk),.wout(w60_124));
	PE pe60_125(.x(x125),.w(w60_124),.acc(r60_124),.res(r60_125),.clk(clk),.wout(w60_125));
	PE pe60_126(.x(x126),.w(w60_125),.acc(r60_125),.res(r60_126),.clk(clk),.wout(w60_126));
	PE pe60_127(.x(x127),.w(w60_126),.acc(r60_126),.res(result60),.clk(clk),.wout(weight60));

	PE pe61_0(.x(x0),.w(w61),.acc(32'h0),.res(r61_0),.clk(clk),.wout(w61_0));
	PE pe61_1(.x(x1),.w(w61_0),.acc(r61_0),.res(r61_1),.clk(clk),.wout(w61_1));
	PE pe61_2(.x(x2),.w(w61_1),.acc(r61_1),.res(r61_2),.clk(clk),.wout(w61_2));
	PE pe61_3(.x(x3),.w(w61_2),.acc(r61_2),.res(r61_3),.clk(clk),.wout(w61_3));
	PE pe61_4(.x(x4),.w(w61_3),.acc(r61_3),.res(r61_4),.clk(clk),.wout(w61_4));
	PE pe61_5(.x(x5),.w(w61_4),.acc(r61_4),.res(r61_5),.clk(clk),.wout(w61_5));
	PE pe61_6(.x(x6),.w(w61_5),.acc(r61_5),.res(r61_6),.clk(clk),.wout(w61_6));
	PE pe61_7(.x(x7),.w(w61_6),.acc(r61_6),.res(r61_7),.clk(clk),.wout(w61_7));
	PE pe61_8(.x(x8),.w(w61_7),.acc(r61_7),.res(r61_8),.clk(clk),.wout(w61_8));
	PE pe61_9(.x(x9),.w(w61_8),.acc(r61_8),.res(r61_9),.clk(clk),.wout(w61_9));
	PE pe61_10(.x(x10),.w(w61_9),.acc(r61_9),.res(r61_10),.clk(clk),.wout(w61_10));
	PE pe61_11(.x(x11),.w(w61_10),.acc(r61_10),.res(r61_11),.clk(clk),.wout(w61_11));
	PE pe61_12(.x(x12),.w(w61_11),.acc(r61_11),.res(r61_12),.clk(clk),.wout(w61_12));
	PE pe61_13(.x(x13),.w(w61_12),.acc(r61_12),.res(r61_13),.clk(clk),.wout(w61_13));
	PE pe61_14(.x(x14),.w(w61_13),.acc(r61_13),.res(r61_14),.clk(clk),.wout(w61_14));
	PE pe61_15(.x(x15),.w(w61_14),.acc(r61_14),.res(r61_15),.clk(clk),.wout(w61_15));
	PE pe61_16(.x(x16),.w(w61_15),.acc(r61_15),.res(r61_16),.clk(clk),.wout(w61_16));
	PE pe61_17(.x(x17),.w(w61_16),.acc(r61_16),.res(r61_17),.clk(clk),.wout(w61_17));
	PE pe61_18(.x(x18),.w(w61_17),.acc(r61_17),.res(r61_18),.clk(clk),.wout(w61_18));
	PE pe61_19(.x(x19),.w(w61_18),.acc(r61_18),.res(r61_19),.clk(clk),.wout(w61_19));
	PE pe61_20(.x(x20),.w(w61_19),.acc(r61_19),.res(r61_20),.clk(clk),.wout(w61_20));
	PE pe61_21(.x(x21),.w(w61_20),.acc(r61_20),.res(r61_21),.clk(clk),.wout(w61_21));
	PE pe61_22(.x(x22),.w(w61_21),.acc(r61_21),.res(r61_22),.clk(clk),.wout(w61_22));
	PE pe61_23(.x(x23),.w(w61_22),.acc(r61_22),.res(r61_23),.clk(clk),.wout(w61_23));
	PE pe61_24(.x(x24),.w(w61_23),.acc(r61_23),.res(r61_24),.clk(clk),.wout(w61_24));
	PE pe61_25(.x(x25),.w(w61_24),.acc(r61_24),.res(r61_25),.clk(clk),.wout(w61_25));
	PE pe61_26(.x(x26),.w(w61_25),.acc(r61_25),.res(r61_26),.clk(clk),.wout(w61_26));
	PE pe61_27(.x(x27),.w(w61_26),.acc(r61_26),.res(r61_27),.clk(clk),.wout(w61_27));
	PE pe61_28(.x(x28),.w(w61_27),.acc(r61_27),.res(r61_28),.clk(clk),.wout(w61_28));
	PE pe61_29(.x(x29),.w(w61_28),.acc(r61_28),.res(r61_29),.clk(clk),.wout(w61_29));
	PE pe61_30(.x(x30),.w(w61_29),.acc(r61_29),.res(r61_30),.clk(clk),.wout(w61_30));
	PE pe61_31(.x(x31),.w(w61_30),.acc(r61_30),.res(r61_31),.clk(clk),.wout(w61_31));
	PE pe61_32(.x(x32),.w(w61_31),.acc(r61_31),.res(r61_32),.clk(clk),.wout(w61_32));
	PE pe61_33(.x(x33),.w(w61_32),.acc(r61_32),.res(r61_33),.clk(clk),.wout(w61_33));
	PE pe61_34(.x(x34),.w(w61_33),.acc(r61_33),.res(r61_34),.clk(clk),.wout(w61_34));
	PE pe61_35(.x(x35),.w(w61_34),.acc(r61_34),.res(r61_35),.clk(clk),.wout(w61_35));
	PE pe61_36(.x(x36),.w(w61_35),.acc(r61_35),.res(r61_36),.clk(clk),.wout(w61_36));
	PE pe61_37(.x(x37),.w(w61_36),.acc(r61_36),.res(r61_37),.clk(clk),.wout(w61_37));
	PE pe61_38(.x(x38),.w(w61_37),.acc(r61_37),.res(r61_38),.clk(clk),.wout(w61_38));
	PE pe61_39(.x(x39),.w(w61_38),.acc(r61_38),.res(r61_39),.clk(clk),.wout(w61_39));
	PE pe61_40(.x(x40),.w(w61_39),.acc(r61_39),.res(r61_40),.clk(clk),.wout(w61_40));
	PE pe61_41(.x(x41),.w(w61_40),.acc(r61_40),.res(r61_41),.clk(clk),.wout(w61_41));
	PE pe61_42(.x(x42),.w(w61_41),.acc(r61_41),.res(r61_42),.clk(clk),.wout(w61_42));
	PE pe61_43(.x(x43),.w(w61_42),.acc(r61_42),.res(r61_43),.clk(clk),.wout(w61_43));
	PE pe61_44(.x(x44),.w(w61_43),.acc(r61_43),.res(r61_44),.clk(clk),.wout(w61_44));
	PE pe61_45(.x(x45),.w(w61_44),.acc(r61_44),.res(r61_45),.clk(clk),.wout(w61_45));
	PE pe61_46(.x(x46),.w(w61_45),.acc(r61_45),.res(r61_46),.clk(clk),.wout(w61_46));
	PE pe61_47(.x(x47),.w(w61_46),.acc(r61_46),.res(r61_47),.clk(clk),.wout(w61_47));
	PE pe61_48(.x(x48),.w(w61_47),.acc(r61_47),.res(r61_48),.clk(clk),.wout(w61_48));
	PE pe61_49(.x(x49),.w(w61_48),.acc(r61_48),.res(r61_49),.clk(clk),.wout(w61_49));
	PE pe61_50(.x(x50),.w(w61_49),.acc(r61_49),.res(r61_50),.clk(clk),.wout(w61_50));
	PE pe61_51(.x(x51),.w(w61_50),.acc(r61_50),.res(r61_51),.clk(clk),.wout(w61_51));
	PE pe61_52(.x(x52),.w(w61_51),.acc(r61_51),.res(r61_52),.clk(clk),.wout(w61_52));
	PE pe61_53(.x(x53),.w(w61_52),.acc(r61_52),.res(r61_53),.clk(clk),.wout(w61_53));
	PE pe61_54(.x(x54),.w(w61_53),.acc(r61_53),.res(r61_54),.clk(clk),.wout(w61_54));
	PE pe61_55(.x(x55),.w(w61_54),.acc(r61_54),.res(r61_55),.clk(clk),.wout(w61_55));
	PE pe61_56(.x(x56),.w(w61_55),.acc(r61_55),.res(r61_56),.clk(clk),.wout(w61_56));
	PE pe61_57(.x(x57),.w(w61_56),.acc(r61_56),.res(r61_57),.clk(clk),.wout(w61_57));
	PE pe61_58(.x(x58),.w(w61_57),.acc(r61_57),.res(r61_58),.clk(clk),.wout(w61_58));
	PE pe61_59(.x(x59),.w(w61_58),.acc(r61_58),.res(r61_59),.clk(clk),.wout(w61_59));
	PE pe61_60(.x(x60),.w(w61_59),.acc(r61_59),.res(r61_60),.clk(clk),.wout(w61_60));
	PE pe61_61(.x(x61),.w(w61_60),.acc(r61_60),.res(r61_61),.clk(clk),.wout(w61_61));
	PE pe61_62(.x(x62),.w(w61_61),.acc(r61_61),.res(r61_62),.clk(clk),.wout(w61_62));
	PE pe61_63(.x(x63),.w(w61_62),.acc(r61_62),.res(r61_63),.clk(clk),.wout(w61_63));
	PE pe61_64(.x(x64),.w(w61_63),.acc(r61_63),.res(r61_64),.clk(clk),.wout(w61_64));
	PE pe61_65(.x(x65),.w(w61_64),.acc(r61_64),.res(r61_65),.clk(clk),.wout(w61_65));
	PE pe61_66(.x(x66),.w(w61_65),.acc(r61_65),.res(r61_66),.clk(clk),.wout(w61_66));
	PE pe61_67(.x(x67),.w(w61_66),.acc(r61_66),.res(r61_67),.clk(clk),.wout(w61_67));
	PE pe61_68(.x(x68),.w(w61_67),.acc(r61_67),.res(r61_68),.clk(clk),.wout(w61_68));
	PE pe61_69(.x(x69),.w(w61_68),.acc(r61_68),.res(r61_69),.clk(clk),.wout(w61_69));
	PE pe61_70(.x(x70),.w(w61_69),.acc(r61_69),.res(r61_70),.clk(clk),.wout(w61_70));
	PE pe61_71(.x(x71),.w(w61_70),.acc(r61_70),.res(r61_71),.clk(clk),.wout(w61_71));
	PE pe61_72(.x(x72),.w(w61_71),.acc(r61_71),.res(r61_72),.clk(clk),.wout(w61_72));
	PE pe61_73(.x(x73),.w(w61_72),.acc(r61_72),.res(r61_73),.clk(clk),.wout(w61_73));
	PE pe61_74(.x(x74),.w(w61_73),.acc(r61_73),.res(r61_74),.clk(clk),.wout(w61_74));
	PE pe61_75(.x(x75),.w(w61_74),.acc(r61_74),.res(r61_75),.clk(clk),.wout(w61_75));
	PE pe61_76(.x(x76),.w(w61_75),.acc(r61_75),.res(r61_76),.clk(clk),.wout(w61_76));
	PE pe61_77(.x(x77),.w(w61_76),.acc(r61_76),.res(r61_77),.clk(clk),.wout(w61_77));
	PE pe61_78(.x(x78),.w(w61_77),.acc(r61_77),.res(r61_78),.clk(clk),.wout(w61_78));
	PE pe61_79(.x(x79),.w(w61_78),.acc(r61_78),.res(r61_79),.clk(clk),.wout(w61_79));
	PE pe61_80(.x(x80),.w(w61_79),.acc(r61_79),.res(r61_80),.clk(clk),.wout(w61_80));
	PE pe61_81(.x(x81),.w(w61_80),.acc(r61_80),.res(r61_81),.clk(clk),.wout(w61_81));
	PE pe61_82(.x(x82),.w(w61_81),.acc(r61_81),.res(r61_82),.clk(clk),.wout(w61_82));
	PE pe61_83(.x(x83),.w(w61_82),.acc(r61_82),.res(r61_83),.clk(clk),.wout(w61_83));
	PE pe61_84(.x(x84),.w(w61_83),.acc(r61_83),.res(r61_84),.clk(clk),.wout(w61_84));
	PE pe61_85(.x(x85),.w(w61_84),.acc(r61_84),.res(r61_85),.clk(clk),.wout(w61_85));
	PE pe61_86(.x(x86),.w(w61_85),.acc(r61_85),.res(r61_86),.clk(clk),.wout(w61_86));
	PE pe61_87(.x(x87),.w(w61_86),.acc(r61_86),.res(r61_87),.clk(clk),.wout(w61_87));
	PE pe61_88(.x(x88),.w(w61_87),.acc(r61_87),.res(r61_88),.clk(clk),.wout(w61_88));
	PE pe61_89(.x(x89),.w(w61_88),.acc(r61_88),.res(r61_89),.clk(clk),.wout(w61_89));
	PE pe61_90(.x(x90),.w(w61_89),.acc(r61_89),.res(r61_90),.clk(clk),.wout(w61_90));
	PE pe61_91(.x(x91),.w(w61_90),.acc(r61_90),.res(r61_91),.clk(clk),.wout(w61_91));
	PE pe61_92(.x(x92),.w(w61_91),.acc(r61_91),.res(r61_92),.clk(clk),.wout(w61_92));
	PE pe61_93(.x(x93),.w(w61_92),.acc(r61_92),.res(r61_93),.clk(clk),.wout(w61_93));
	PE pe61_94(.x(x94),.w(w61_93),.acc(r61_93),.res(r61_94),.clk(clk),.wout(w61_94));
	PE pe61_95(.x(x95),.w(w61_94),.acc(r61_94),.res(r61_95),.clk(clk),.wout(w61_95));
	PE pe61_96(.x(x96),.w(w61_95),.acc(r61_95),.res(r61_96),.clk(clk),.wout(w61_96));
	PE pe61_97(.x(x97),.w(w61_96),.acc(r61_96),.res(r61_97),.clk(clk),.wout(w61_97));
	PE pe61_98(.x(x98),.w(w61_97),.acc(r61_97),.res(r61_98),.clk(clk),.wout(w61_98));
	PE pe61_99(.x(x99),.w(w61_98),.acc(r61_98),.res(r61_99),.clk(clk),.wout(w61_99));
	PE pe61_100(.x(x100),.w(w61_99),.acc(r61_99),.res(r61_100),.clk(clk),.wout(w61_100));
	PE pe61_101(.x(x101),.w(w61_100),.acc(r61_100),.res(r61_101),.clk(clk),.wout(w61_101));
	PE pe61_102(.x(x102),.w(w61_101),.acc(r61_101),.res(r61_102),.clk(clk),.wout(w61_102));
	PE pe61_103(.x(x103),.w(w61_102),.acc(r61_102),.res(r61_103),.clk(clk),.wout(w61_103));
	PE pe61_104(.x(x104),.w(w61_103),.acc(r61_103),.res(r61_104),.clk(clk),.wout(w61_104));
	PE pe61_105(.x(x105),.w(w61_104),.acc(r61_104),.res(r61_105),.clk(clk),.wout(w61_105));
	PE pe61_106(.x(x106),.w(w61_105),.acc(r61_105),.res(r61_106),.clk(clk),.wout(w61_106));
	PE pe61_107(.x(x107),.w(w61_106),.acc(r61_106),.res(r61_107),.clk(clk),.wout(w61_107));
	PE pe61_108(.x(x108),.w(w61_107),.acc(r61_107),.res(r61_108),.clk(clk),.wout(w61_108));
	PE pe61_109(.x(x109),.w(w61_108),.acc(r61_108),.res(r61_109),.clk(clk),.wout(w61_109));
	PE pe61_110(.x(x110),.w(w61_109),.acc(r61_109),.res(r61_110),.clk(clk),.wout(w61_110));
	PE pe61_111(.x(x111),.w(w61_110),.acc(r61_110),.res(r61_111),.clk(clk),.wout(w61_111));
	PE pe61_112(.x(x112),.w(w61_111),.acc(r61_111),.res(r61_112),.clk(clk),.wout(w61_112));
	PE pe61_113(.x(x113),.w(w61_112),.acc(r61_112),.res(r61_113),.clk(clk),.wout(w61_113));
	PE pe61_114(.x(x114),.w(w61_113),.acc(r61_113),.res(r61_114),.clk(clk),.wout(w61_114));
	PE pe61_115(.x(x115),.w(w61_114),.acc(r61_114),.res(r61_115),.clk(clk),.wout(w61_115));
	PE pe61_116(.x(x116),.w(w61_115),.acc(r61_115),.res(r61_116),.clk(clk),.wout(w61_116));
	PE pe61_117(.x(x117),.w(w61_116),.acc(r61_116),.res(r61_117),.clk(clk),.wout(w61_117));
	PE pe61_118(.x(x118),.w(w61_117),.acc(r61_117),.res(r61_118),.clk(clk),.wout(w61_118));
	PE pe61_119(.x(x119),.w(w61_118),.acc(r61_118),.res(r61_119),.clk(clk),.wout(w61_119));
	PE pe61_120(.x(x120),.w(w61_119),.acc(r61_119),.res(r61_120),.clk(clk),.wout(w61_120));
	PE pe61_121(.x(x121),.w(w61_120),.acc(r61_120),.res(r61_121),.clk(clk),.wout(w61_121));
	PE pe61_122(.x(x122),.w(w61_121),.acc(r61_121),.res(r61_122),.clk(clk),.wout(w61_122));
	PE pe61_123(.x(x123),.w(w61_122),.acc(r61_122),.res(r61_123),.clk(clk),.wout(w61_123));
	PE pe61_124(.x(x124),.w(w61_123),.acc(r61_123),.res(r61_124),.clk(clk),.wout(w61_124));
	PE pe61_125(.x(x125),.w(w61_124),.acc(r61_124),.res(r61_125),.clk(clk),.wout(w61_125));
	PE pe61_126(.x(x126),.w(w61_125),.acc(r61_125),.res(r61_126),.clk(clk),.wout(w61_126));
	PE pe61_127(.x(x127),.w(w61_126),.acc(r61_126),.res(result61),.clk(clk),.wout(weight61));

	PE pe62_0(.x(x0),.w(w62),.acc(32'h0),.res(r62_0),.clk(clk),.wout(w62_0));
	PE pe62_1(.x(x1),.w(w62_0),.acc(r62_0),.res(r62_1),.clk(clk),.wout(w62_1));
	PE pe62_2(.x(x2),.w(w62_1),.acc(r62_1),.res(r62_2),.clk(clk),.wout(w62_2));
	PE pe62_3(.x(x3),.w(w62_2),.acc(r62_2),.res(r62_3),.clk(clk),.wout(w62_3));
	PE pe62_4(.x(x4),.w(w62_3),.acc(r62_3),.res(r62_4),.clk(clk),.wout(w62_4));
	PE pe62_5(.x(x5),.w(w62_4),.acc(r62_4),.res(r62_5),.clk(clk),.wout(w62_5));
	PE pe62_6(.x(x6),.w(w62_5),.acc(r62_5),.res(r62_6),.clk(clk),.wout(w62_6));
	PE pe62_7(.x(x7),.w(w62_6),.acc(r62_6),.res(r62_7),.clk(clk),.wout(w62_7));
	PE pe62_8(.x(x8),.w(w62_7),.acc(r62_7),.res(r62_8),.clk(clk),.wout(w62_8));
	PE pe62_9(.x(x9),.w(w62_8),.acc(r62_8),.res(r62_9),.clk(clk),.wout(w62_9));
	PE pe62_10(.x(x10),.w(w62_9),.acc(r62_9),.res(r62_10),.clk(clk),.wout(w62_10));
	PE pe62_11(.x(x11),.w(w62_10),.acc(r62_10),.res(r62_11),.clk(clk),.wout(w62_11));
	PE pe62_12(.x(x12),.w(w62_11),.acc(r62_11),.res(r62_12),.clk(clk),.wout(w62_12));
	PE pe62_13(.x(x13),.w(w62_12),.acc(r62_12),.res(r62_13),.clk(clk),.wout(w62_13));
	PE pe62_14(.x(x14),.w(w62_13),.acc(r62_13),.res(r62_14),.clk(clk),.wout(w62_14));
	PE pe62_15(.x(x15),.w(w62_14),.acc(r62_14),.res(r62_15),.clk(clk),.wout(w62_15));
	PE pe62_16(.x(x16),.w(w62_15),.acc(r62_15),.res(r62_16),.clk(clk),.wout(w62_16));
	PE pe62_17(.x(x17),.w(w62_16),.acc(r62_16),.res(r62_17),.clk(clk),.wout(w62_17));
	PE pe62_18(.x(x18),.w(w62_17),.acc(r62_17),.res(r62_18),.clk(clk),.wout(w62_18));
	PE pe62_19(.x(x19),.w(w62_18),.acc(r62_18),.res(r62_19),.clk(clk),.wout(w62_19));
	PE pe62_20(.x(x20),.w(w62_19),.acc(r62_19),.res(r62_20),.clk(clk),.wout(w62_20));
	PE pe62_21(.x(x21),.w(w62_20),.acc(r62_20),.res(r62_21),.clk(clk),.wout(w62_21));
	PE pe62_22(.x(x22),.w(w62_21),.acc(r62_21),.res(r62_22),.clk(clk),.wout(w62_22));
	PE pe62_23(.x(x23),.w(w62_22),.acc(r62_22),.res(r62_23),.clk(clk),.wout(w62_23));
	PE pe62_24(.x(x24),.w(w62_23),.acc(r62_23),.res(r62_24),.clk(clk),.wout(w62_24));
	PE pe62_25(.x(x25),.w(w62_24),.acc(r62_24),.res(r62_25),.clk(clk),.wout(w62_25));
	PE pe62_26(.x(x26),.w(w62_25),.acc(r62_25),.res(r62_26),.clk(clk),.wout(w62_26));
	PE pe62_27(.x(x27),.w(w62_26),.acc(r62_26),.res(r62_27),.clk(clk),.wout(w62_27));
	PE pe62_28(.x(x28),.w(w62_27),.acc(r62_27),.res(r62_28),.clk(clk),.wout(w62_28));
	PE pe62_29(.x(x29),.w(w62_28),.acc(r62_28),.res(r62_29),.clk(clk),.wout(w62_29));
	PE pe62_30(.x(x30),.w(w62_29),.acc(r62_29),.res(r62_30),.clk(clk),.wout(w62_30));
	PE pe62_31(.x(x31),.w(w62_30),.acc(r62_30),.res(r62_31),.clk(clk),.wout(w62_31));
	PE pe62_32(.x(x32),.w(w62_31),.acc(r62_31),.res(r62_32),.clk(clk),.wout(w62_32));
	PE pe62_33(.x(x33),.w(w62_32),.acc(r62_32),.res(r62_33),.clk(clk),.wout(w62_33));
	PE pe62_34(.x(x34),.w(w62_33),.acc(r62_33),.res(r62_34),.clk(clk),.wout(w62_34));
	PE pe62_35(.x(x35),.w(w62_34),.acc(r62_34),.res(r62_35),.clk(clk),.wout(w62_35));
	PE pe62_36(.x(x36),.w(w62_35),.acc(r62_35),.res(r62_36),.clk(clk),.wout(w62_36));
	PE pe62_37(.x(x37),.w(w62_36),.acc(r62_36),.res(r62_37),.clk(clk),.wout(w62_37));
	PE pe62_38(.x(x38),.w(w62_37),.acc(r62_37),.res(r62_38),.clk(clk),.wout(w62_38));
	PE pe62_39(.x(x39),.w(w62_38),.acc(r62_38),.res(r62_39),.clk(clk),.wout(w62_39));
	PE pe62_40(.x(x40),.w(w62_39),.acc(r62_39),.res(r62_40),.clk(clk),.wout(w62_40));
	PE pe62_41(.x(x41),.w(w62_40),.acc(r62_40),.res(r62_41),.clk(clk),.wout(w62_41));
	PE pe62_42(.x(x42),.w(w62_41),.acc(r62_41),.res(r62_42),.clk(clk),.wout(w62_42));
	PE pe62_43(.x(x43),.w(w62_42),.acc(r62_42),.res(r62_43),.clk(clk),.wout(w62_43));
	PE pe62_44(.x(x44),.w(w62_43),.acc(r62_43),.res(r62_44),.clk(clk),.wout(w62_44));
	PE pe62_45(.x(x45),.w(w62_44),.acc(r62_44),.res(r62_45),.clk(clk),.wout(w62_45));
	PE pe62_46(.x(x46),.w(w62_45),.acc(r62_45),.res(r62_46),.clk(clk),.wout(w62_46));
	PE pe62_47(.x(x47),.w(w62_46),.acc(r62_46),.res(r62_47),.clk(clk),.wout(w62_47));
	PE pe62_48(.x(x48),.w(w62_47),.acc(r62_47),.res(r62_48),.clk(clk),.wout(w62_48));
	PE pe62_49(.x(x49),.w(w62_48),.acc(r62_48),.res(r62_49),.clk(clk),.wout(w62_49));
	PE pe62_50(.x(x50),.w(w62_49),.acc(r62_49),.res(r62_50),.clk(clk),.wout(w62_50));
	PE pe62_51(.x(x51),.w(w62_50),.acc(r62_50),.res(r62_51),.clk(clk),.wout(w62_51));
	PE pe62_52(.x(x52),.w(w62_51),.acc(r62_51),.res(r62_52),.clk(clk),.wout(w62_52));
	PE pe62_53(.x(x53),.w(w62_52),.acc(r62_52),.res(r62_53),.clk(clk),.wout(w62_53));
	PE pe62_54(.x(x54),.w(w62_53),.acc(r62_53),.res(r62_54),.clk(clk),.wout(w62_54));
	PE pe62_55(.x(x55),.w(w62_54),.acc(r62_54),.res(r62_55),.clk(clk),.wout(w62_55));
	PE pe62_56(.x(x56),.w(w62_55),.acc(r62_55),.res(r62_56),.clk(clk),.wout(w62_56));
	PE pe62_57(.x(x57),.w(w62_56),.acc(r62_56),.res(r62_57),.clk(clk),.wout(w62_57));
	PE pe62_58(.x(x58),.w(w62_57),.acc(r62_57),.res(r62_58),.clk(clk),.wout(w62_58));
	PE pe62_59(.x(x59),.w(w62_58),.acc(r62_58),.res(r62_59),.clk(clk),.wout(w62_59));
	PE pe62_60(.x(x60),.w(w62_59),.acc(r62_59),.res(r62_60),.clk(clk),.wout(w62_60));
	PE pe62_61(.x(x61),.w(w62_60),.acc(r62_60),.res(r62_61),.clk(clk),.wout(w62_61));
	PE pe62_62(.x(x62),.w(w62_61),.acc(r62_61),.res(r62_62),.clk(clk),.wout(w62_62));
	PE pe62_63(.x(x63),.w(w62_62),.acc(r62_62),.res(r62_63),.clk(clk),.wout(w62_63));
	PE pe62_64(.x(x64),.w(w62_63),.acc(r62_63),.res(r62_64),.clk(clk),.wout(w62_64));
	PE pe62_65(.x(x65),.w(w62_64),.acc(r62_64),.res(r62_65),.clk(clk),.wout(w62_65));
	PE pe62_66(.x(x66),.w(w62_65),.acc(r62_65),.res(r62_66),.clk(clk),.wout(w62_66));
	PE pe62_67(.x(x67),.w(w62_66),.acc(r62_66),.res(r62_67),.clk(clk),.wout(w62_67));
	PE pe62_68(.x(x68),.w(w62_67),.acc(r62_67),.res(r62_68),.clk(clk),.wout(w62_68));
	PE pe62_69(.x(x69),.w(w62_68),.acc(r62_68),.res(r62_69),.clk(clk),.wout(w62_69));
	PE pe62_70(.x(x70),.w(w62_69),.acc(r62_69),.res(r62_70),.clk(clk),.wout(w62_70));
	PE pe62_71(.x(x71),.w(w62_70),.acc(r62_70),.res(r62_71),.clk(clk),.wout(w62_71));
	PE pe62_72(.x(x72),.w(w62_71),.acc(r62_71),.res(r62_72),.clk(clk),.wout(w62_72));
	PE pe62_73(.x(x73),.w(w62_72),.acc(r62_72),.res(r62_73),.clk(clk),.wout(w62_73));
	PE pe62_74(.x(x74),.w(w62_73),.acc(r62_73),.res(r62_74),.clk(clk),.wout(w62_74));
	PE pe62_75(.x(x75),.w(w62_74),.acc(r62_74),.res(r62_75),.clk(clk),.wout(w62_75));
	PE pe62_76(.x(x76),.w(w62_75),.acc(r62_75),.res(r62_76),.clk(clk),.wout(w62_76));
	PE pe62_77(.x(x77),.w(w62_76),.acc(r62_76),.res(r62_77),.clk(clk),.wout(w62_77));
	PE pe62_78(.x(x78),.w(w62_77),.acc(r62_77),.res(r62_78),.clk(clk),.wout(w62_78));
	PE pe62_79(.x(x79),.w(w62_78),.acc(r62_78),.res(r62_79),.clk(clk),.wout(w62_79));
	PE pe62_80(.x(x80),.w(w62_79),.acc(r62_79),.res(r62_80),.clk(clk),.wout(w62_80));
	PE pe62_81(.x(x81),.w(w62_80),.acc(r62_80),.res(r62_81),.clk(clk),.wout(w62_81));
	PE pe62_82(.x(x82),.w(w62_81),.acc(r62_81),.res(r62_82),.clk(clk),.wout(w62_82));
	PE pe62_83(.x(x83),.w(w62_82),.acc(r62_82),.res(r62_83),.clk(clk),.wout(w62_83));
	PE pe62_84(.x(x84),.w(w62_83),.acc(r62_83),.res(r62_84),.clk(clk),.wout(w62_84));
	PE pe62_85(.x(x85),.w(w62_84),.acc(r62_84),.res(r62_85),.clk(clk),.wout(w62_85));
	PE pe62_86(.x(x86),.w(w62_85),.acc(r62_85),.res(r62_86),.clk(clk),.wout(w62_86));
	PE pe62_87(.x(x87),.w(w62_86),.acc(r62_86),.res(r62_87),.clk(clk),.wout(w62_87));
	PE pe62_88(.x(x88),.w(w62_87),.acc(r62_87),.res(r62_88),.clk(clk),.wout(w62_88));
	PE pe62_89(.x(x89),.w(w62_88),.acc(r62_88),.res(r62_89),.clk(clk),.wout(w62_89));
	PE pe62_90(.x(x90),.w(w62_89),.acc(r62_89),.res(r62_90),.clk(clk),.wout(w62_90));
	PE pe62_91(.x(x91),.w(w62_90),.acc(r62_90),.res(r62_91),.clk(clk),.wout(w62_91));
	PE pe62_92(.x(x92),.w(w62_91),.acc(r62_91),.res(r62_92),.clk(clk),.wout(w62_92));
	PE pe62_93(.x(x93),.w(w62_92),.acc(r62_92),.res(r62_93),.clk(clk),.wout(w62_93));
	PE pe62_94(.x(x94),.w(w62_93),.acc(r62_93),.res(r62_94),.clk(clk),.wout(w62_94));
	PE pe62_95(.x(x95),.w(w62_94),.acc(r62_94),.res(r62_95),.clk(clk),.wout(w62_95));
	PE pe62_96(.x(x96),.w(w62_95),.acc(r62_95),.res(r62_96),.clk(clk),.wout(w62_96));
	PE pe62_97(.x(x97),.w(w62_96),.acc(r62_96),.res(r62_97),.clk(clk),.wout(w62_97));
	PE pe62_98(.x(x98),.w(w62_97),.acc(r62_97),.res(r62_98),.clk(clk),.wout(w62_98));
	PE pe62_99(.x(x99),.w(w62_98),.acc(r62_98),.res(r62_99),.clk(clk),.wout(w62_99));
	PE pe62_100(.x(x100),.w(w62_99),.acc(r62_99),.res(r62_100),.clk(clk),.wout(w62_100));
	PE pe62_101(.x(x101),.w(w62_100),.acc(r62_100),.res(r62_101),.clk(clk),.wout(w62_101));
	PE pe62_102(.x(x102),.w(w62_101),.acc(r62_101),.res(r62_102),.clk(clk),.wout(w62_102));
	PE pe62_103(.x(x103),.w(w62_102),.acc(r62_102),.res(r62_103),.clk(clk),.wout(w62_103));
	PE pe62_104(.x(x104),.w(w62_103),.acc(r62_103),.res(r62_104),.clk(clk),.wout(w62_104));
	PE pe62_105(.x(x105),.w(w62_104),.acc(r62_104),.res(r62_105),.clk(clk),.wout(w62_105));
	PE pe62_106(.x(x106),.w(w62_105),.acc(r62_105),.res(r62_106),.clk(clk),.wout(w62_106));
	PE pe62_107(.x(x107),.w(w62_106),.acc(r62_106),.res(r62_107),.clk(clk),.wout(w62_107));
	PE pe62_108(.x(x108),.w(w62_107),.acc(r62_107),.res(r62_108),.clk(clk),.wout(w62_108));
	PE pe62_109(.x(x109),.w(w62_108),.acc(r62_108),.res(r62_109),.clk(clk),.wout(w62_109));
	PE pe62_110(.x(x110),.w(w62_109),.acc(r62_109),.res(r62_110),.clk(clk),.wout(w62_110));
	PE pe62_111(.x(x111),.w(w62_110),.acc(r62_110),.res(r62_111),.clk(clk),.wout(w62_111));
	PE pe62_112(.x(x112),.w(w62_111),.acc(r62_111),.res(r62_112),.clk(clk),.wout(w62_112));
	PE pe62_113(.x(x113),.w(w62_112),.acc(r62_112),.res(r62_113),.clk(clk),.wout(w62_113));
	PE pe62_114(.x(x114),.w(w62_113),.acc(r62_113),.res(r62_114),.clk(clk),.wout(w62_114));
	PE pe62_115(.x(x115),.w(w62_114),.acc(r62_114),.res(r62_115),.clk(clk),.wout(w62_115));
	PE pe62_116(.x(x116),.w(w62_115),.acc(r62_115),.res(r62_116),.clk(clk),.wout(w62_116));
	PE pe62_117(.x(x117),.w(w62_116),.acc(r62_116),.res(r62_117),.clk(clk),.wout(w62_117));
	PE pe62_118(.x(x118),.w(w62_117),.acc(r62_117),.res(r62_118),.clk(clk),.wout(w62_118));
	PE pe62_119(.x(x119),.w(w62_118),.acc(r62_118),.res(r62_119),.clk(clk),.wout(w62_119));
	PE pe62_120(.x(x120),.w(w62_119),.acc(r62_119),.res(r62_120),.clk(clk),.wout(w62_120));
	PE pe62_121(.x(x121),.w(w62_120),.acc(r62_120),.res(r62_121),.clk(clk),.wout(w62_121));
	PE pe62_122(.x(x122),.w(w62_121),.acc(r62_121),.res(r62_122),.clk(clk),.wout(w62_122));
	PE pe62_123(.x(x123),.w(w62_122),.acc(r62_122),.res(r62_123),.clk(clk),.wout(w62_123));
	PE pe62_124(.x(x124),.w(w62_123),.acc(r62_123),.res(r62_124),.clk(clk),.wout(w62_124));
	PE pe62_125(.x(x125),.w(w62_124),.acc(r62_124),.res(r62_125),.clk(clk),.wout(w62_125));
	PE pe62_126(.x(x126),.w(w62_125),.acc(r62_125),.res(r62_126),.clk(clk),.wout(w62_126));
	PE pe62_127(.x(x127),.w(w62_126),.acc(r62_126),.res(result62),.clk(clk),.wout(weight62));

	PE pe63_0(.x(x0),.w(w63),.acc(32'h0),.res(r63_0),.clk(clk),.wout(w63_0));
	PE pe63_1(.x(x1),.w(w63_0),.acc(r63_0),.res(r63_1),.clk(clk),.wout(w63_1));
	PE pe63_2(.x(x2),.w(w63_1),.acc(r63_1),.res(r63_2),.clk(clk),.wout(w63_2));
	PE pe63_3(.x(x3),.w(w63_2),.acc(r63_2),.res(r63_3),.clk(clk),.wout(w63_3));
	PE pe63_4(.x(x4),.w(w63_3),.acc(r63_3),.res(r63_4),.clk(clk),.wout(w63_4));
	PE pe63_5(.x(x5),.w(w63_4),.acc(r63_4),.res(r63_5),.clk(clk),.wout(w63_5));
	PE pe63_6(.x(x6),.w(w63_5),.acc(r63_5),.res(r63_6),.clk(clk),.wout(w63_6));
	PE pe63_7(.x(x7),.w(w63_6),.acc(r63_6),.res(r63_7),.clk(clk),.wout(w63_7));
	PE pe63_8(.x(x8),.w(w63_7),.acc(r63_7),.res(r63_8),.clk(clk),.wout(w63_8));
	PE pe63_9(.x(x9),.w(w63_8),.acc(r63_8),.res(r63_9),.clk(clk),.wout(w63_9));
	PE pe63_10(.x(x10),.w(w63_9),.acc(r63_9),.res(r63_10),.clk(clk),.wout(w63_10));
	PE pe63_11(.x(x11),.w(w63_10),.acc(r63_10),.res(r63_11),.clk(clk),.wout(w63_11));
	PE pe63_12(.x(x12),.w(w63_11),.acc(r63_11),.res(r63_12),.clk(clk),.wout(w63_12));
	PE pe63_13(.x(x13),.w(w63_12),.acc(r63_12),.res(r63_13),.clk(clk),.wout(w63_13));
	PE pe63_14(.x(x14),.w(w63_13),.acc(r63_13),.res(r63_14),.clk(clk),.wout(w63_14));
	PE pe63_15(.x(x15),.w(w63_14),.acc(r63_14),.res(r63_15),.clk(clk),.wout(w63_15));
	PE pe63_16(.x(x16),.w(w63_15),.acc(r63_15),.res(r63_16),.clk(clk),.wout(w63_16));
	PE pe63_17(.x(x17),.w(w63_16),.acc(r63_16),.res(r63_17),.clk(clk),.wout(w63_17));
	PE pe63_18(.x(x18),.w(w63_17),.acc(r63_17),.res(r63_18),.clk(clk),.wout(w63_18));
	PE pe63_19(.x(x19),.w(w63_18),.acc(r63_18),.res(r63_19),.clk(clk),.wout(w63_19));
	PE pe63_20(.x(x20),.w(w63_19),.acc(r63_19),.res(r63_20),.clk(clk),.wout(w63_20));
	PE pe63_21(.x(x21),.w(w63_20),.acc(r63_20),.res(r63_21),.clk(clk),.wout(w63_21));
	PE pe63_22(.x(x22),.w(w63_21),.acc(r63_21),.res(r63_22),.clk(clk),.wout(w63_22));
	PE pe63_23(.x(x23),.w(w63_22),.acc(r63_22),.res(r63_23),.clk(clk),.wout(w63_23));
	PE pe63_24(.x(x24),.w(w63_23),.acc(r63_23),.res(r63_24),.clk(clk),.wout(w63_24));
	PE pe63_25(.x(x25),.w(w63_24),.acc(r63_24),.res(r63_25),.clk(clk),.wout(w63_25));
	PE pe63_26(.x(x26),.w(w63_25),.acc(r63_25),.res(r63_26),.clk(clk),.wout(w63_26));
	PE pe63_27(.x(x27),.w(w63_26),.acc(r63_26),.res(r63_27),.clk(clk),.wout(w63_27));
	PE pe63_28(.x(x28),.w(w63_27),.acc(r63_27),.res(r63_28),.clk(clk),.wout(w63_28));
	PE pe63_29(.x(x29),.w(w63_28),.acc(r63_28),.res(r63_29),.clk(clk),.wout(w63_29));
	PE pe63_30(.x(x30),.w(w63_29),.acc(r63_29),.res(r63_30),.clk(clk),.wout(w63_30));
	PE pe63_31(.x(x31),.w(w63_30),.acc(r63_30),.res(r63_31),.clk(clk),.wout(w63_31));
	PE pe63_32(.x(x32),.w(w63_31),.acc(r63_31),.res(r63_32),.clk(clk),.wout(w63_32));
	PE pe63_33(.x(x33),.w(w63_32),.acc(r63_32),.res(r63_33),.clk(clk),.wout(w63_33));
	PE pe63_34(.x(x34),.w(w63_33),.acc(r63_33),.res(r63_34),.clk(clk),.wout(w63_34));
	PE pe63_35(.x(x35),.w(w63_34),.acc(r63_34),.res(r63_35),.clk(clk),.wout(w63_35));
	PE pe63_36(.x(x36),.w(w63_35),.acc(r63_35),.res(r63_36),.clk(clk),.wout(w63_36));
	PE pe63_37(.x(x37),.w(w63_36),.acc(r63_36),.res(r63_37),.clk(clk),.wout(w63_37));
	PE pe63_38(.x(x38),.w(w63_37),.acc(r63_37),.res(r63_38),.clk(clk),.wout(w63_38));
	PE pe63_39(.x(x39),.w(w63_38),.acc(r63_38),.res(r63_39),.clk(clk),.wout(w63_39));
	PE pe63_40(.x(x40),.w(w63_39),.acc(r63_39),.res(r63_40),.clk(clk),.wout(w63_40));
	PE pe63_41(.x(x41),.w(w63_40),.acc(r63_40),.res(r63_41),.clk(clk),.wout(w63_41));
	PE pe63_42(.x(x42),.w(w63_41),.acc(r63_41),.res(r63_42),.clk(clk),.wout(w63_42));
	PE pe63_43(.x(x43),.w(w63_42),.acc(r63_42),.res(r63_43),.clk(clk),.wout(w63_43));
	PE pe63_44(.x(x44),.w(w63_43),.acc(r63_43),.res(r63_44),.clk(clk),.wout(w63_44));
	PE pe63_45(.x(x45),.w(w63_44),.acc(r63_44),.res(r63_45),.clk(clk),.wout(w63_45));
	PE pe63_46(.x(x46),.w(w63_45),.acc(r63_45),.res(r63_46),.clk(clk),.wout(w63_46));
	PE pe63_47(.x(x47),.w(w63_46),.acc(r63_46),.res(r63_47),.clk(clk),.wout(w63_47));
	PE pe63_48(.x(x48),.w(w63_47),.acc(r63_47),.res(r63_48),.clk(clk),.wout(w63_48));
	PE pe63_49(.x(x49),.w(w63_48),.acc(r63_48),.res(r63_49),.clk(clk),.wout(w63_49));
	PE pe63_50(.x(x50),.w(w63_49),.acc(r63_49),.res(r63_50),.clk(clk),.wout(w63_50));
	PE pe63_51(.x(x51),.w(w63_50),.acc(r63_50),.res(r63_51),.clk(clk),.wout(w63_51));
	PE pe63_52(.x(x52),.w(w63_51),.acc(r63_51),.res(r63_52),.clk(clk),.wout(w63_52));
	PE pe63_53(.x(x53),.w(w63_52),.acc(r63_52),.res(r63_53),.clk(clk),.wout(w63_53));
	PE pe63_54(.x(x54),.w(w63_53),.acc(r63_53),.res(r63_54),.clk(clk),.wout(w63_54));
	PE pe63_55(.x(x55),.w(w63_54),.acc(r63_54),.res(r63_55),.clk(clk),.wout(w63_55));
	PE pe63_56(.x(x56),.w(w63_55),.acc(r63_55),.res(r63_56),.clk(clk),.wout(w63_56));
	PE pe63_57(.x(x57),.w(w63_56),.acc(r63_56),.res(r63_57),.clk(clk),.wout(w63_57));
	PE pe63_58(.x(x58),.w(w63_57),.acc(r63_57),.res(r63_58),.clk(clk),.wout(w63_58));
	PE pe63_59(.x(x59),.w(w63_58),.acc(r63_58),.res(r63_59),.clk(clk),.wout(w63_59));
	PE pe63_60(.x(x60),.w(w63_59),.acc(r63_59),.res(r63_60),.clk(clk),.wout(w63_60));
	PE pe63_61(.x(x61),.w(w63_60),.acc(r63_60),.res(r63_61),.clk(clk),.wout(w63_61));
	PE pe63_62(.x(x62),.w(w63_61),.acc(r63_61),.res(r63_62),.clk(clk),.wout(w63_62));
	PE pe63_63(.x(x63),.w(w63_62),.acc(r63_62),.res(r63_63),.clk(clk),.wout(w63_63));
	PE pe63_64(.x(x64),.w(w63_63),.acc(r63_63),.res(r63_64),.clk(clk),.wout(w63_64));
	PE pe63_65(.x(x65),.w(w63_64),.acc(r63_64),.res(r63_65),.clk(clk),.wout(w63_65));
	PE pe63_66(.x(x66),.w(w63_65),.acc(r63_65),.res(r63_66),.clk(clk),.wout(w63_66));
	PE pe63_67(.x(x67),.w(w63_66),.acc(r63_66),.res(r63_67),.clk(clk),.wout(w63_67));
	PE pe63_68(.x(x68),.w(w63_67),.acc(r63_67),.res(r63_68),.clk(clk),.wout(w63_68));
	PE pe63_69(.x(x69),.w(w63_68),.acc(r63_68),.res(r63_69),.clk(clk),.wout(w63_69));
	PE pe63_70(.x(x70),.w(w63_69),.acc(r63_69),.res(r63_70),.clk(clk),.wout(w63_70));
	PE pe63_71(.x(x71),.w(w63_70),.acc(r63_70),.res(r63_71),.clk(clk),.wout(w63_71));
	PE pe63_72(.x(x72),.w(w63_71),.acc(r63_71),.res(r63_72),.clk(clk),.wout(w63_72));
	PE pe63_73(.x(x73),.w(w63_72),.acc(r63_72),.res(r63_73),.clk(clk),.wout(w63_73));
	PE pe63_74(.x(x74),.w(w63_73),.acc(r63_73),.res(r63_74),.clk(clk),.wout(w63_74));
	PE pe63_75(.x(x75),.w(w63_74),.acc(r63_74),.res(r63_75),.clk(clk),.wout(w63_75));
	PE pe63_76(.x(x76),.w(w63_75),.acc(r63_75),.res(r63_76),.clk(clk),.wout(w63_76));
	PE pe63_77(.x(x77),.w(w63_76),.acc(r63_76),.res(r63_77),.clk(clk),.wout(w63_77));
	PE pe63_78(.x(x78),.w(w63_77),.acc(r63_77),.res(r63_78),.clk(clk),.wout(w63_78));
	PE pe63_79(.x(x79),.w(w63_78),.acc(r63_78),.res(r63_79),.clk(clk),.wout(w63_79));
	PE pe63_80(.x(x80),.w(w63_79),.acc(r63_79),.res(r63_80),.clk(clk),.wout(w63_80));
	PE pe63_81(.x(x81),.w(w63_80),.acc(r63_80),.res(r63_81),.clk(clk),.wout(w63_81));
	PE pe63_82(.x(x82),.w(w63_81),.acc(r63_81),.res(r63_82),.clk(clk),.wout(w63_82));
	PE pe63_83(.x(x83),.w(w63_82),.acc(r63_82),.res(r63_83),.clk(clk),.wout(w63_83));
	PE pe63_84(.x(x84),.w(w63_83),.acc(r63_83),.res(r63_84),.clk(clk),.wout(w63_84));
	PE pe63_85(.x(x85),.w(w63_84),.acc(r63_84),.res(r63_85),.clk(clk),.wout(w63_85));
	PE pe63_86(.x(x86),.w(w63_85),.acc(r63_85),.res(r63_86),.clk(clk),.wout(w63_86));
	PE pe63_87(.x(x87),.w(w63_86),.acc(r63_86),.res(r63_87),.clk(clk),.wout(w63_87));
	PE pe63_88(.x(x88),.w(w63_87),.acc(r63_87),.res(r63_88),.clk(clk),.wout(w63_88));
	PE pe63_89(.x(x89),.w(w63_88),.acc(r63_88),.res(r63_89),.clk(clk),.wout(w63_89));
	PE pe63_90(.x(x90),.w(w63_89),.acc(r63_89),.res(r63_90),.clk(clk),.wout(w63_90));
	PE pe63_91(.x(x91),.w(w63_90),.acc(r63_90),.res(r63_91),.clk(clk),.wout(w63_91));
	PE pe63_92(.x(x92),.w(w63_91),.acc(r63_91),.res(r63_92),.clk(clk),.wout(w63_92));
	PE pe63_93(.x(x93),.w(w63_92),.acc(r63_92),.res(r63_93),.clk(clk),.wout(w63_93));
	PE pe63_94(.x(x94),.w(w63_93),.acc(r63_93),.res(r63_94),.clk(clk),.wout(w63_94));
	PE pe63_95(.x(x95),.w(w63_94),.acc(r63_94),.res(r63_95),.clk(clk),.wout(w63_95));
	PE pe63_96(.x(x96),.w(w63_95),.acc(r63_95),.res(r63_96),.clk(clk),.wout(w63_96));
	PE pe63_97(.x(x97),.w(w63_96),.acc(r63_96),.res(r63_97),.clk(clk),.wout(w63_97));
	PE pe63_98(.x(x98),.w(w63_97),.acc(r63_97),.res(r63_98),.clk(clk),.wout(w63_98));
	PE pe63_99(.x(x99),.w(w63_98),.acc(r63_98),.res(r63_99),.clk(clk),.wout(w63_99));
	PE pe63_100(.x(x100),.w(w63_99),.acc(r63_99),.res(r63_100),.clk(clk),.wout(w63_100));
	PE pe63_101(.x(x101),.w(w63_100),.acc(r63_100),.res(r63_101),.clk(clk),.wout(w63_101));
	PE pe63_102(.x(x102),.w(w63_101),.acc(r63_101),.res(r63_102),.clk(clk),.wout(w63_102));
	PE pe63_103(.x(x103),.w(w63_102),.acc(r63_102),.res(r63_103),.clk(clk),.wout(w63_103));
	PE pe63_104(.x(x104),.w(w63_103),.acc(r63_103),.res(r63_104),.clk(clk),.wout(w63_104));
	PE pe63_105(.x(x105),.w(w63_104),.acc(r63_104),.res(r63_105),.clk(clk),.wout(w63_105));
	PE pe63_106(.x(x106),.w(w63_105),.acc(r63_105),.res(r63_106),.clk(clk),.wout(w63_106));
	PE pe63_107(.x(x107),.w(w63_106),.acc(r63_106),.res(r63_107),.clk(clk),.wout(w63_107));
	PE pe63_108(.x(x108),.w(w63_107),.acc(r63_107),.res(r63_108),.clk(clk),.wout(w63_108));
	PE pe63_109(.x(x109),.w(w63_108),.acc(r63_108),.res(r63_109),.clk(clk),.wout(w63_109));
	PE pe63_110(.x(x110),.w(w63_109),.acc(r63_109),.res(r63_110),.clk(clk),.wout(w63_110));
	PE pe63_111(.x(x111),.w(w63_110),.acc(r63_110),.res(r63_111),.clk(clk),.wout(w63_111));
	PE pe63_112(.x(x112),.w(w63_111),.acc(r63_111),.res(r63_112),.clk(clk),.wout(w63_112));
	PE pe63_113(.x(x113),.w(w63_112),.acc(r63_112),.res(r63_113),.clk(clk),.wout(w63_113));
	PE pe63_114(.x(x114),.w(w63_113),.acc(r63_113),.res(r63_114),.clk(clk),.wout(w63_114));
	PE pe63_115(.x(x115),.w(w63_114),.acc(r63_114),.res(r63_115),.clk(clk),.wout(w63_115));
	PE pe63_116(.x(x116),.w(w63_115),.acc(r63_115),.res(r63_116),.clk(clk),.wout(w63_116));
	PE pe63_117(.x(x117),.w(w63_116),.acc(r63_116),.res(r63_117),.clk(clk),.wout(w63_117));
	PE pe63_118(.x(x118),.w(w63_117),.acc(r63_117),.res(r63_118),.clk(clk),.wout(w63_118));
	PE pe63_119(.x(x119),.w(w63_118),.acc(r63_118),.res(r63_119),.clk(clk),.wout(w63_119));
	PE pe63_120(.x(x120),.w(w63_119),.acc(r63_119),.res(r63_120),.clk(clk),.wout(w63_120));
	PE pe63_121(.x(x121),.w(w63_120),.acc(r63_120),.res(r63_121),.clk(clk),.wout(w63_121));
	PE pe63_122(.x(x122),.w(w63_121),.acc(r63_121),.res(r63_122),.clk(clk),.wout(w63_122));
	PE pe63_123(.x(x123),.w(w63_122),.acc(r63_122),.res(r63_123),.clk(clk),.wout(w63_123));
	PE pe63_124(.x(x124),.w(w63_123),.acc(r63_123),.res(r63_124),.clk(clk),.wout(w63_124));
	PE pe63_125(.x(x125),.w(w63_124),.acc(r63_124),.res(r63_125),.clk(clk),.wout(w63_125));
	PE pe63_126(.x(x126),.w(w63_125),.acc(r63_125),.res(r63_126),.clk(clk),.wout(w63_126));
	PE pe63_127(.x(x127),.w(w63_126),.acc(r63_126),.res(result63),.clk(clk),.wout(weight63));

	PE pe64_0(.x(x0),.w(w64),.acc(32'h0),.res(r64_0),.clk(clk),.wout(w64_0));
	PE pe64_1(.x(x1),.w(w64_0),.acc(r64_0),.res(r64_1),.clk(clk),.wout(w64_1));
	PE pe64_2(.x(x2),.w(w64_1),.acc(r64_1),.res(r64_2),.clk(clk),.wout(w64_2));
	PE pe64_3(.x(x3),.w(w64_2),.acc(r64_2),.res(r64_3),.clk(clk),.wout(w64_3));
	PE pe64_4(.x(x4),.w(w64_3),.acc(r64_3),.res(r64_4),.clk(clk),.wout(w64_4));
	PE pe64_5(.x(x5),.w(w64_4),.acc(r64_4),.res(r64_5),.clk(clk),.wout(w64_5));
	PE pe64_6(.x(x6),.w(w64_5),.acc(r64_5),.res(r64_6),.clk(clk),.wout(w64_6));
	PE pe64_7(.x(x7),.w(w64_6),.acc(r64_6),.res(r64_7),.clk(clk),.wout(w64_7));
	PE pe64_8(.x(x8),.w(w64_7),.acc(r64_7),.res(r64_8),.clk(clk),.wout(w64_8));
	PE pe64_9(.x(x9),.w(w64_8),.acc(r64_8),.res(r64_9),.clk(clk),.wout(w64_9));
	PE pe64_10(.x(x10),.w(w64_9),.acc(r64_9),.res(r64_10),.clk(clk),.wout(w64_10));
	PE pe64_11(.x(x11),.w(w64_10),.acc(r64_10),.res(r64_11),.clk(clk),.wout(w64_11));
	PE pe64_12(.x(x12),.w(w64_11),.acc(r64_11),.res(r64_12),.clk(clk),.wout(w64_12));
	PE pe64_13(.x(x13),.w(w64_12),.acc(r64_12),.res(r64_13),.clk(clk),.wout(w64_13));
	PE pe64_14(.x(x14),.w(w64_13),.acc(r64_13),.res(r64_14),.clk(clk),.wout(w64_14));
	PE pe64_15(.x(x15),.w(w64_14),.acc(r64_14),.res(r64_15),.clk(clk),.wout(w64_15));
	PE pe64_16(.x(x16),.w(w64_15),.acc(r64_15),.res(r64_16),.clk(clk),.wout(w64_16));
	PE pe64_17(.x(x17),.w(w64_16),.acc(r64_16),.res(r64_17),.clk(clk),.wout(w64_17));
	PE pe64_18(.x(x18),.w(w64_17),.acc(r64_17),.res(r64_18),.clk(clk),.wout(w64_18));
	PE pe64_19(.x(x19),.w(w64_18),.acc(r64_18),.res(r64_19),.clk(clk),.wout(w64_19));
	PE pe64_20(.x(x20),.w(w64_19),.acc(r64_19),.res(r64_20),.clk(clk),.wout(w64_20));
	PE pe64_21(.x(x21),.w(w64_20),.acc(r64_20),.res(r64_21),.clk(clk),.wout(w64_21));
	PE pe64_22(.x(x22),.w(w64_21),.acc(r64_21),.res(r64_22),.clk(clk),.wout(w64_22));
	PE pe64_23(.x(x23),.w(w64_22),.acc(r64_22),.res(r64_23),.clk(clk),.wout(w64_23));
	PE pe64_24(.x(x24),.w(w64_23),.acc(r64_23),.res(r64_24),.clk(clk),.wout(w64_24));
	PE pe64_25(.x(x25),.w(w64_24),.acc(r64_24),.res(r64_25),.clk(clk),.wout(w64_25));
	PE pe64_26(.x(x26),.w(w64_25),.acc(r64_25),.res(r64_26),.clk(clk),.wout(w64_26));
	PE pe64_27(.x(x27),.w(w64_26),.acc(r64_26),.res(r64_27),.clk(clk),.wout(w64_27));
	PE pe64_28(.x(x28),.w(w64_27),.acc(r64_27),.res(r64_28),.clk(clk),.wout(w64_28));
	PE pe64_29(.x(x29),.w(w64_28),.acc(r64_28),.res(r64_29),.clk(clk),.wout(w64_29));
	PE pe64_30(.x(x30),.w(w64_29),.acc(r64_29),.res(r64_30),.clk(clk),.wout(w64_30));
	PE pe64_31(.x(x31),.w(w64_30),.acc(r64_30),.res(r64_31),.clk(clk),.wout(w64_31));
	PE pe64_32(.x(x32),.w(w64_31),.acc(r64_31),.res(r64_32),.clk(clk),.wout(w64_32));
	PE pe64_33(.x(x33),.w(w64_32),.acc(r64_32),.res(r64_33),.clk(clk),.wout(w64_33));
	PE pe64_34(.x(x34),.w(w64_33),.acc(r64_33),.res(r64_34),.clk(clk),.wout(w64_34));
	PE pe64_35(.x(x35),.w(w64_34),.acc(r64_34),.res(r64_35),.clk(clk),.wout(w64_35));
	PE pe64_36(.x(x36),.w(w64_35),.acc(r64_35),.res(r64_36),.clk(clk),.wout(w64_36));
	PE pe64_37(.x(x37),.w(w64_36),.acc(r64_36),.res(r64_37),.clk(clk),.wout(w64_37));
	PE pe64_38(.x(x38),.w(w64_37),.acc(r64_37),.res(r64_38),.clk(clk),.wout(w64_38));
	PE pe64_39(.x(x39),.w(w64_38),.acc(r64_38),.res(r64_39),.clk(clk),.wout(w64_39));
	PE pe64_40(.x(x40),.w(w64_39),.acc(r64_39),.res(r64_40),.clk(clk),.wout(w64_40));
	PE pe64_41(.x(x41),.w(w64_40),.acc(r64_40),.res(r64_41),.clk(clk),.wout(w64_41));
	PE pe64_42(.x(x42),.w(w64_41),.acc(r64_41),.res(r64_42),.clk(clk),.wout(w64_42));
	PE pe64_43(.x(x43),.w(w64_42),.acc(r64_42),.res(r64_43),.clk(clk),.wout(w64_43));
	PE pe64_44(.x(x44),.w(w64_43),.acc(r64_43),.res(r64_44),.clk(clk),.wout(w64_44));
	PE pe64_45(.x(x45),.w(w64_44),.acc(r64_44),.res(r64_45),.clk(clk),.wout(w64_45));
	PE pe64_46(.x(x46),.w(w64_45),.acc(r64_45),.res(r64_46),.clk(clk),.wout(w64_46));
	PE pe64_47(.x(x47),.w(w64_46),.acc(r64_46),.res(r64_47),.clk(clk),.wout(w64_47));
	PE pe64_48(.x(x48),.w(w64_47),.acc(r64_47),.res(r64_48),.clk(clk),.wout(w64_48));
	PE pe64_49(.x(x49),.w(w64_48),.acc(r64_48),.res(r64_49),.clk(clk),.wout(w64_49));
	PE pe64_50(.x(x50),.w(w64_49),.acc(r64_49),.res(r64_50),.clk(clk),.wout(w64_50));
	PE pe64_51(.x(x51),.w(w64_50),.acc(r64_50),.res(r64_51),.clk(clk),.wout(w64_51));
	PE pe64_52(.x(x52),.w(w64_51),.acc(r64_51),.res(r64_52),.clk(clk),.wout(w64_52));
	PE pe64_53(.x(x53),.w(w64_52),.acc(r64_52),.res(r64_53),.clk(clk),.wout(w64_53));
	PE pe64_54(.x(x54),.w(w64_53),.acc(r64_53),.res(r64_54),.clk(clk),.wout(w64_54));
	PE pe64_55(.x(x55),.w(w64_54),.acc(r64_54),.res(r64_55),.clk(clk),.wout(w64_55));
	PE pe64_56(.x(x56),.w(w64_55),.acc(r64_55),.res(r64_56),.clk(clk),.wout(w64_56));
	PE pe64_57(.x(x57),.w(w64_56),.acc(r64_56),.res(r64_57),.clk(clk),.wout(w64_57));
	PE pe64_58(.x(x58),.w(w64_57),.acc(r64_57),.res(r64_58),.clk(clk),.wout(w64_58));
	PE pe64_59(.x(x59),.w(w64_58),.acc(r64_58),.res(r64_59),.clk(clk),.wout(w64_59));
	PE pe64_60(.x(x60),.w(w64_59),.acc(r64_59),.res(r64_60),.clk(clk),.wout(w64_60));
	PE pe64_61(.x(x61),.w(w64_60),.acc(r64_60),.res(r64_61),.clk(clk),.wout(w64_61));
	PE pe64_62(.x(x62),.w(w64_61),.acc(r64_61),.res(r64_62),.clk(clk),.wout(w64_62));
	PE pe64_63(.x(x63),.w(w64_62),.acc(r64_62),.res(r64_63),.clk(clk),.wout(w64_63));
	PE pe64_64(.x(x64),.w(w64_63),.acc(r64_63),.res(r64_64),.clk(clk),.wout(w64_64));
	PE pe64_65(.x(x65),.w(w64_64),.acc(r64_64),.res(r64_65),.clk(clk),.wout(w64_65));
	PE pe64_66(.x(x66),.w(w64_65),.acc(r64_65),.res(r64_66),.clk(clk),.wout(w64_66));
	PE pe64_67(.x(x67),.w(w64_66),.acc(r64_66),.res(r64_67),.clk(clk),.wout(w64_67));
	PE pe64_68(.x(x68),.w(w64_67),.acc(r64_67),.res(r64_68),.clk(clk),.wout(w64_68));
	PE pe64_69(.x(x69),.w(w64_68),.acc(r64_68),.res(r64_69),.clk(clk),.wout(w64_69));
	PE pe64_70(.x(x70),.w(w64_69),.acc(r64_69),.res(r64_70),.clk(clk),.wout(w64_70));
	PE pe64_71(.x(x71),.w(w64_70),.acc(r64_70),.res(r64_71),.clk(clk),.wout(w64_71));
	PE pe64_72(.x(x72),.w(w64_71),.acc(r64_71),.res(r64_72),.clk(clk),.wout(w64_72));
	PE pe64_73(.x(x73),.w(w64_72),.acc(r64_72),.res(r64_73),.clk(clk),.wout(w64_73));
	PE pe64_74(.x(x74),.w(w64_73),.acc(r64_73),.res(r64_74),.clk(clk),.wout(w64_74));
	PE pe64_75(.x(x75),.w(w64_74),.acc(r64_74),.res(r64_75),.clk(clk),.wout(w64_75));
	PE pe64_76(.x(x76),.w(w64_75),.acc(r64_75),.res(r64_76),.clk(clk),.wout(w64_76));
	PE pe64_77(.x(x77),.w(w64_76),.acc(r64_76),.res(r64_77),.clk(clk),.wout(w64_77));
	PE pe64_78(.x(x78),.w(w64_77),.acc(r64_77),.res(r64_78),.clk(clk),.wout(w64_78));
	PE pe64_79(.x(x79),.w(w64_78),.acc(r64_78),.res(r64_79),.clk(clk),.wout(w64_79));
	PE pe64_80(.x(x80),.w(w64_79),.acc(r64_79),.res(r64_80),.clk(clk),.wout(w64_80));
	PE pe64_81(.x(x81),.w(w64_80),.acc(r64_80),.res(r64_81),.clk(clk),.wout(w64_81));
	PE pe64_82(.x(x82),.w(w64_81),.acc(r64_81),.res(r64_82),.clk(clk),.wout(w64_82));
	PE pe64_83(.x(x83),.w(w64_82),.acc(r64_82),.res(r64_83),.clk(clk),.wout(w64_83));
	PE pe64_84(.x(x84),.w(w64_83),.acc(r64_83),.res(r64_84),.clk(clk),.wout(w64_84));
	PE pe64_85(.x(x85),.w(w64_84),.acc(r64_84),.res(r64_85),.clk(clk),.wout(w64_85));
	PE pe64_86(.x(x86),.w(w64_85),.acc(r64_85),.res(r64_86),.clk(clk),.wout(w64_86));
	PE pe64_87(.x(x87),.w(w64_86),.acc(r64_86),.res(r64_87),.clk(clk),.wout(w64_87));
	PE pe64_88(.x(x88),.w(w64_87),.acc(r64_87),.res(r64_88),.clk(clk),.wout(w64_88));
	PE pe64_89(.x(x89),.w(w64_88),.acc(r64_88),.res(r64_89),.clk(clk),.wout(w64_89));
	PE pe64_90(.x(x90),.w(w64_89),.acc(r64_89),.res(r64_90),.clk(clk),.wout(w64_90));
	PE pe64_91(.x(x91),.w(w64_90),.acc(r64_90),.res(r64_91),.clk(clk),.wout(w64_91));
	PE pe64_92(.x(x92),.w(w64_91),.acc(r64_91),.res(r64_92),.clk(clk),.wout(w64_92));
	PE pe64_93(.x(x93),.w(w64_92),.acc(r64_92),.res(r64_93),.clk(clk),.wout(w64_93));
	PE pe64_94(.x(x94),.w(w64_93),.acc(r64_93),.res(r64_94),.clk(clk),.wout(w64_94));
	PE pe64_95(.x(x95),.w(w64_94),.acc(r64_94),.res(r64_95),.clk(clk),.wout(w64_95));
	PE pe64_96(.x(x96),.w(w64_95),.acc(r64_95),.res(r64_96),.clk(clk),.wout(w64_96));
	PE pe64_97(.x(x97),.w(w64_96),.acc(r64_96),.res(r64_97),.clk(clk),.wout(w64_97));
	PE pe64_98(.x(x98),.w(w64_97),.acc(r64_97),.res(r64_98),.clk(clk),.wout(w64_98));
	PE pe64_99(.x(x99),.w(w64_98),.acc(r64_98),.res(r64_99),.clk(clk),.wout(w64_99));
	PE pe64_100(.x(x100),.w(w64_99),.acc(r64_99),.res(r64_100),.clk(clk),.wout(w64_100));
	PE pe64_101(.x(x101),.w(w64_100),.acc(r64_100),.res(r64_101),.clk(clk),.wout(w64_101));
	PE pe64_102(.x(x102),.w(w64_101),.acc(r64_101),.res(r64_102),.clk(clk),.wout(w64_102));
	PE pe64_103(.x(x103),.w(w64_102),.acc(r64_102),.res(r64_103),.clk(clk),.wout(w64_103));
	PE pe64_104(.x(x104),.w(w64_103),.acc(r64_103),.res(r64_104),.clk(clk),.wout(w64_104));
	PE pe64_105(.x(x105),.w(w64_104),.acc(r64_104),.res(r64_105),.clk(clk),.wout(w64_105));
	PE pe64_106(.x(x106),.w(w64_105),.acc(r64_105),.res(r64_106),.clk(clk),.wout(w64_106));
	PE pe64_107(.x(x107),.w(w64_106),.acc(r64_106),.res(r64_107),.clk(clk),.wout(w64_107));
	PE pe64_108(.x(x108),.w(w64_107),.acc(r64_107),.res(r64_108),.clk(clk),.wout(w64_108));
	PE pe64_109(.x(x109),.w(w64_108),.acc(r64_108),.res(r64_109),.clk(clk),.wout(w64_109));
	PE pe64_110(.x(x110),.w(w64_109),.acc(r64_109),.res(r64_110),.clk(clk),.wout(w64_110));
	PE pe64_111(.x(x111),.w(w64_110),.acc(r64_110),.res(r64_111),.clk(clk),.wout(w64_111));
	PE pe64_112(.x(x112),.w(w64_111),.acc(r64_111),.res(r64_112),.clk(clk),.wout(w64_112));
	PE pe64_113(.x(x113),.w(w64_112),.acc(r64_112),.res(r64_113),.clk(clk),.wout(w64_113));
	PE pe64_114(.x(x114),.w(w64_113),.acc(r64_113),.res(r64_114),.clk(clk),.wout(w64_114));
	PE pe64_115(.x(x115),.w(w64_114),.acc(r64_114),.res(r64_115),.clk(clk),.wout(w64_115));
	PE pe64_116(.x(x116),.w(w64_115),.acc(r64_115),.res(r64_116),.clk(clk),.wout(w64_116));
	PE pe64_117(.x(x117),.w(w64_116),.acc(r64_116),.res(r64_117),.clk(clk),.wout(w64_117));
	PE pe64_118(.x(x118),.w(w64_117),.acc(r64_117),.res(r64_118),.clk(clk),.wout(w64_118));
	PE pe64_119(.x(x119),.w(w64_118),.acc(r64_118),.res(r64_119),.clk(clk),.wout(w64_119));
	PE pe64_120(.x(x120),.w(w64_119),.acc(r64_119),.res(r64_120),.clk(clk),.wout(w64_120));
	PE pe64_121(.x(x121),.w(w64_120),.acc(r64_120),.res(r64_121),.clk(clk),.wout(w64_121));
	PE pe64_122(.x(x122),.w(w64_121),.acc(r64_121),.res(r64_122),.clk(clk),.wout(w64_122));
	PE pe64_123(.x(x123),.w(w64_122),.acc(r64_122),.res(r64_123),.clk(clk),.wout(w64_123));
	PE pe64_124(.x(x124),.w(w64_123),.acc(r64_123),.res(r64_124),.clk(clk),.wout(w64_124));
	PE pe64_125(.x(x125),.w(w64_124),.acc(r64_124),.res(r64_125),.clk(clk),.wout(w64_125));
	PE pe64_126(.x(x126),.w(w64_125),.acc(r64_125),.res(r64_126),.clk(clk),.wout(w64_126));
	PE pe64_127(.x(x127),.w(w64_126),.acc(r64_126),.res(result64),.clk(clk),.wout(weight64));

	PE pe65_0(.x(x0),.w(w65),.acc(32'h0),.res(r65_0),.clk(clk),.wout(w65_0));
	PE pe65_1(.x(x1),.w(w65_0),.acc(r65_0),.res(r65_1),.clk(clk),.wout(w65_1));
	PE pe65_2(.x(x2),.w(w65_1),.acc(r65_1),.res(r65_2),.clk(clk),.wout(w65_2));
	PE pe65_3(.x(x3),.w(w65_2),.acc(r65_2),.res(r65_3),.clk(clk),.wout(w65_3));
	PE pe65_4(.x(x4),.w(w65_3),.acc(r65_3),.res(r65_4),.clk(clk),.wout(w65_4));
	PE pe65_5(.x(x5),.w(w65_4),.acc(r65_4),.res(r65_5),.clk(clk),.wout(w65_5));
	PE pe65_6(.x(x6),.w(w65_5),.acc(r65_5),.res(r65_6),.clk(clk),.wout(w65_6));
	PE pe65_7(.x(x7),.w(w65_6),.acc(r65_6),.res(r65_7),.clk(clk),.wout(w65_7));
	PE pe65_8(.x(x8),.w(w65_7),.acc(r65_7),.res(r65_8),.clk(clk),.wout(w65_8));
	PE pe65_9(.x(x9),.w(w65_8),.acc(r65_8),.res(r65_9),.clk(clk),.wout(w65_9));
	PE pe65_10(.x(x10),.w(w65_9),.acc(r65_9),.res(r65_10),.clk(clk),.wout(w65_10));
	PE pe65_11(.x(x11),.w(w65_10),.acc(r65_10),.res(r65_11),.clk(clk),.wout(w65_11));
	PE pe65_12(.x(x12),.w(w65_11),.acc(r65_11),.res(r65_12),.clk(clk),.wout(w65_12));
	PE pe65_13(.x(x13),.w(w65_12),.acc(r65_12),.res(r65_13),.clk(clk),.wout(w65_13));
	PE pe65_14(.x(x14),.w(w65_13),.acc(r65_13),.res(r65_14),.clk(clk),.wout(w65_14));
	PE pe65_15(.x(x15),.w(w65_14),.acc(r65_14),.res(r65_15),.clk(clk),.wout(w65_15));
	PE pe65_16(.x(x16),.w(w65_15),.acc(r65_15),.res(r65_16),.clk(clk),.wout(w65_16));
	PE pe65_17(.x(x17),.w(w65_16),.acc(r65_16),.res(r65_17),.clk(clk),.wout(w65_17));
	PE pe65_18(.x(x18),.w(w65_17),.acc(r65_17),.res(r65_18),.clk(clk),.wout(w65_18));
	PE pe65_19(.x(x19),.w(w65_18),.acc(r65_18),.res(r65_19),.clk(clk),.wout(w65_19));
	PE pe65_20(.x(x20),.w(w65_19),.acc(r65_19),.res(r65_20),.clk(clk),.wout(w65_20));
	PE pe65_21(.x(x21),.w(w65_20),.acc(r65_20),.res(r65_21),.clk(clk),.wout(w65_21));
	PE pe65_22(.x(x22),.w(w65_21),.acc(r65_21),.res(r65_22),.clk(clk),.wout(w65_22));
	PE pe65_23(.x(x23),.w(w65_22),.acc(r65_22),.res(r65_23),.clk(clk),.wout(w65_23));
	PE pe65_24(.x(x24),.w(w65_23),.acc(r65_23),.res(r65_24),.clk(clk),.wout(w65_24));
	PE pe65_25(.x(x25),.w(w65_24),.acc(r65_24),.res(r65_25),.clk(clk),.wout(w65_25));
	PE pe65_26(.x(x26),.w(w65_25),.acc(r65_25),.res(r65_26),.clk(clk),.wout(w65_26));
	PE pe65_27(.x(x27),.w(w65_26),.acc(r65_26),.res(r65_27),.clk(clk),.wout(w65_27));
	PE pe65_28(.x(x28),.w(w65_27),.acc(r65_27),.res(r65_28),.clk(clk),.wout(w65_28));
	PE pe65_29(.x(x29),.w(w65_28),.acc(r65_28),.res(r65_29),.clk(clk),.wout(w65_29));
	PE pe65_30(.x(x30),.w(w65_29),.acc(r65_29),.res(r65_30),.clk(clk),.wout(w65_30));
	PE pe65_31(.x(x31),.w(w65_30),.acc(r65_30),.res(r65_31),.clk(clk),.wout(w65_31));
	PE pe65_32(.x(x32),.w(w65_31),.acc(r65_31),.res(r65_32),.clk(clk),.wout(w65_32));
	PE pe65_33(.x(x33),.w(w65_32),.acc(r65_32),.res(r65_33),.clk(clk),.wout(w65_33));
	PE pe65_34(.x(x34),.w(w65_33),.acc(r65_33),.res(r65_34),.clk(clk),.wout(w65_34));
	PE pe65_35(.x(x35),.w(w65_34),.acc(r65_34),.res(r65_35),.clk(clk),.wout(w65_35));
	PE pe65_36(.x(x36),.w(w65_35),.acc(r65_35),.res(r65_36),.clk(clk),.wout(w65_36));
	PE pe65_37(.x(x37),.w(w65_36),.acc(r65_36),.res(r65_37),.clk(clk),.wout(w65_37));
	PE pe65_38(.x(x38),.w(w65_37),.acc(r65_37),.res(r65_38),.clk(clk),.wout(w65_38));
	PE pe65_39(.x(x39),.w(w65_38),.acc(r65_38),.res(r65_39),.clk(clk),.wout(w65_39));
	PE pe65_40(.x(x40),.w(w65_39),.acc(r65_39),.res(r65_40),.clk(clk),.wout(w65_40));
	PE pe65_41(.x(x41),.w(w65_40),.acc(r65_40),.res(r65_41),.clk(clk),.wout(w65_41));
	PE pe65_42(.x(x42),.w(w65_41),.acc(r65_41),.res(r65_42),.clk(clk),.wout(w65_42));
	PE pe65_43(.x(x43),.w(w65_42),.acc(r65_42),.res(r65_43),.clk(clk),.wout(w65_43));
	PE pe65_44(.x(x44),.w(w65_43),.acc(r65_43),.res(r65_44),.clk(clk),.wout(w65_44));
	PE pe65_45(.x(x45),.w(w65_44),.acc(r65_44),.res(r65_45),.clk(clk),.wout(w65_45));
	PE pe65_46(.x(x46),.w(w65_45),.acc(r65_45),.res(r65_46),.clk(clk),.wout(w65_46));
	PE pe65_47(.x(x47),.w(w65_46),.acc(r65_46),.res(r65_47),.clk(clk),.wout(w65_47));
	PE pe65_48(.x(x48),.w(w65_47),.acc(r65_47),.res(r65_48),.clk(clk),.wout(w65_48));
	PE pe65_49(.x(x49),.w(w65_48),.acc(r65_48),.res(r65_49),.clk(clk),.wout(w65_49));
	PE pe65_50(.x(x50),.w(w65_49),.acc(r65_49),.res(r65_50),.clk(clk),.wout(w65_50));
	PE pe65_51(.x(x51),.w(w65_50),.acc(r65_50),.res(r65_51),.clk(clk),.wout(w65_51));
	PE pe65_52(.x(x52),.w(w65_51),.acc(r65_51),.res(r65_52),.clk(clk),.wout(w65_52));
	PE pe65_53(.x(x53),.w(w65_52),.acc(r65_52),.res(r65_53),.clk(clk),.wout(w65_53));
	PE pe65_54(.x(x54),.w(w65_53),.acc(r65_53),.res(r65_54),.clk(clk),.wout(w65_54));
	PE pe65_55(.x(x55),.w(w65_54),.acc(r65_54),.res(r65_55),.clk(clk),.wout(w65_55));
	PE pe65_56(.x(x56),.w(w65_55),.acc(r65_55),.res(r65_56),.clk(clk),.wout(w65_56));
	PE pe65_57(.x(x57),.w(w65_56),.acc(r65_56),.res(r65_57),.clk(clk),.wout(w65_57));
	PE pe65_58(.x(x58),.w(w65_57),.acc(r65_57),.res(r65_58),.clk(clk),.wout(w65_58));
	PE pe65_59(.x(x59),.w(w65_58),.acc(r65_58),.res(r65_59),.clk(clk),.wout(w65_59));
	PE pe65_60(.x(x60),.w(w65_59),.acc(r65_59),.res(r65_60),.clk(clk),.wout(w65_60));
	PE pe65_61(.x(x61),.w(w65_60),.acc(r65_60),.res(r65_61),.clk(clk),.wout(w65_61));
	PE pe65_62(.x(x62),.w(w65_61),.acc(r65_61),.res(r65_62),.clk(clk),.wout(w65_62));
	PE pe65_63(.x(x63),.w(w65_62),.acc(r65_62),.res(r65_63),.clk(clk),.wout(w65_63));
	PE pe65_64(.x(x64),.w(w65_63),.acc(r65_63),.res(r65_64),.clk(clk),.wout(w65_64));
	PE pe65_65(.x(x65),.w(w65_64),.acc(r65_64),.res(r65_65),.clk(clk),.wout(w65_65));
	PE pe65_66(.x(x66),.w(w65_65),.acc(r65_65),.res(r65_66),.clk(clk),.wout(w65_66));
	PE pe65_67(.x(x67),.w(w65_66),.acc(r65_66),.res(r65_67),.clk(clk),.wout(w65_67));
	PE pe65_68(.x(x68),.w(w65_67),.acc(r65_67),.res(r65_68),.clk(clk),.wout(w65_68));
	PE pe65_69(.x(x69),.w(w65_68),.acc(r65_68),.res(r65_69),.clk(clk),.wout(w65_69));
	PE pe65_70(.x(x70),.w(w65_69),.acc(r65_69),.res(r65_70),.clk(clk),.wout(w65_70));
	PE pe65_71(.x(x71),.w(w65_70),.acc(r65_70),.res(r65_71),.clk(clk),.wout(w65_71));
	PE pe65_72(.x(x72),.w(w65_71),.acc(r65_71),.res(r65_72),.clk(clk),.wout(w65_72));
	PE pe65_73(.x(x73),.w(w65_72),.acc(r65_72),.res(r65_73),.clk(clk),.wout(w65_73));
	PE pe65_74(.x(x74),.w(w65_73),.acc(r65_73),.res(r65_74),.clk(clk),.wout(w65_74));
	PE pe65_75(.x(x75),.w(w65_74),.acc(r65_74),.res(r65_75),.clk(clk),.wout(w65_75));
	PE pe65_76(.x(x76),.w(w65_75),.acc(r65_75),.res(r65_76),.clk(clk),.wout(w65_76));
	PE pe65_77(.x(x77),.w(w65_76),.acc(r65_76),.res(r65_77),.clk(clk),.wout(w65_77));
	PE pe65_78(.x(x78),.w(w65_77),.acc(r65_77),.res(r65_78),.clk(clk),.wout(w65_78));
	PE pe65_79(.x(x79),.w(w65_78),.acc(r65_78),.res(r65_79),.clk(clk),.wout(w65_79));
	PE pe65_80(.x(x80),.w(w65_79),.acc(r65_79),.res(r65_80),.clk(clk),.wout(w65_80));
	PE pe65_81(.x(x81),.w(w65_80),.acc(r65_80),.res(r65_81),.clk(clk),.wout(w65_81));
	PE pe65_82(.x(x82),.w(w65_81),.acc(r65_81),.res(r65_82),.clk(clk),.wout(w65_82));
	PE pe65_83(.x(x83),.w(w65_82),.acc(r65_82),.res(r65_83),.clk(clk),.wout(w65_83));
	PE pe65_84(.x(x84),.w(w65_83),.acc(r65_83),.res(r65_84),.clk(clk),.wout(w65_84));
	PE pe65_85(.x(x85),.w(w65_84),.acc(r65_84),.res(r65_85),.clk(clk),.wout(w65_85));
	PE pe65_86(.x(x86),.w(w65_85),.acc(r65_85),.res(r65_86),.clk(clk),.wout(w65_86));
	PE pe65_87(.x(x87),.w(w65_86),.acc(r65_86),.res(r65_87),.clk(clk),.wout(w65_87));
	PE pe65_88(.x(x88),.w(w65_87),.acc(r65_87),.res(r65_88),.clk(clk),.wout(w65_88));
	PE pe65_89(.x(x89),.w(w65_88),.acc(r65_88),.res(r65_89),.clk(clk),.wout(w65_89));
	PE pe65_90(.x(x90),.w(w65_89),.acc(r65_89),.res(r65_90),.clk(clk),.wout(w65_90));
	PE pe65_91(.x(x91),.w(w65_90),.acc(r65_90),.res(r65_91),.clk(clk),.wout(w65_91));
	PE pe65_92(.x(x92),.w(w65_91),.acc(r65_91),.res(r65_92),.clk(clk),.wout(w65_92));
	PE pe65_93(.x(x93),.w(w65_92),.acc(r65_92),.res(r65_93),.clk(clk),.wout(w65_93));
	PE pe65_94(.x(x94),.w(w65_93),.acc(r65_93),.res(r65_94),.clk(clk),.wout(w65_94));
	PE pe65_95(.x(x95),.w(w65_94),.acc(r65_94),.res(r65_95),.clk(clk),.wout(w65_95));
	PE pe65_96(.x(x96),.w(w65_95),.acc(r65_95),.res(r65_96),.clk(clk),.wout(w65_96));
	PE pe65_97(.x(x97),.w(w65_96),.acc(r65_96),.res(r65_97),.clk(clk),.wout(w65_97));
	PE pe65_98(.x(x98),.w(w65_97),.acc(r65_97),.res(r65_98),.clk(clk),.wout(w65_98));
	PE pe65_99(.x(x99),.w(w65_98),.acc(r65_98),.res(r65_99),.clk(clk),.wout(w65_99));
	PE pe65_100(.x(x100),.w(w65_99),.acc(r65_99),.res(r65_100),.clk(clk),.wout(w65_100));
	PE pe65_101(.x(x101),.w(w65_100),.acc(r65_100),.res(r65_101),.clk(clk),.wout(w65_101));
	PE pe65_102(.x(x102),.w(w65_101),.acc(r65_101),.res(r65_102),.clk(clk),.wout(w65_102));
	PE pe65_103(.x(x103),.w(w65_102),.acc(r65_102),.res(r65_103),.clk(clk),.wout(w65_103));
	PE pe65_104(.x(x104),.w(w65_103),.acc(r65_103),.res(r65_104),.clk(clk),.wout(w65_104));
	PE pe65_105(.x(x105),.w(w65_104),.acc(r65_104),.res(r65_105),.clk(clk),.wout(w65_105));
	PE pe65_106(.x(x106),.w(w65_105),.acc(r65_105),.res(r65_106),.clk(clk),.wout(w65_106));
	PE pe65_107(.x(x107),.w(w65_106),.acc(r65_106),.res(r65_107),.clk(clk),.wout(w65_107));
	PE pe65_108(.x(x108),.w(w65_107),.acc(r65_107),.res(r65_108),.clk(clk),.wout(w65_108));
	PE pe65_109(.x(x109),.w(w65_108),.acc(r65_108),.res(r65_109),.clk(clk),.wout(w65_109));
	PE pe65_110(.x(x110),.w(w65_109),.acc(r65_109),.res(r65_110),.clk(clk),.wout(w65_110));
	PE pe65_111(.x(x111),.w(w65_110),.acc(r65_110),.res(r65_111),.clk(clk),.wout(w65_111));
	PE pe65_112(.x(x112),.w(w65_111),.acc(r65_111),.res(r65_112),.clk(clk),.wout(w65_112));
	PE pe65_113(.x(x113),.w(w65_112),.acc(r65_112),.res(r65_113),.clk(clk),.wout(w65_113));
	PE pe65_114(.x(x114),.w(w65_113),.acc(r65_113),.res(r65_114),.clk(clk),.wout(w65_114));
	PE pe65_115(.x(x115),.w(w65_114),.acc(r65_114),.res(r65_115),.clk(clk),.wout(w65_115));
	PE pe65_116(.x(x116),.w(w65_115),.acc(r65_115),.res(r65_116),.clk(clk),.wout(w65_116));
	PE pe65_117(.x(x117),.w(w65_116),.acc(r65_116),.res(r65_117),.clk(clk),.wout(w65_117));
	PE pe65_118(.x(x118),.w(w65_117),.acc(r65_117),.res(r65_118),.clk(clk),.wout(w65_118));
	PE pe65_119(.x(x119),.w(w65_118),.acc(r65_118),.res(r65_119),.clk(clk),.wout(w65_119));
	PE pe65_120(.x(x120),.w(w65_119),.acc(r65_119),.res(r65_120),.clk(clk),.wout(w65_120));
	PE pe65_121(.x(x121),.w(w65_120),.acc(r65_120),.res(r65_121),.clk(clk),.wout(w65_121));
	PE pe65_122(.x(x122),.w(w65_121),.acc(r65_121),.res(r65_122),.clk(clk),.wout(w65_122));
	PE pe65_123(.x(x123),.w(w65_122),.acc(r65_122),.res(r65_123),.clk(clk),.wout(w65_123));
	PE pe65_124(.x(x124),.w(w65_123),.acc(r65_123),.res(r65_124),.clk(clk),.wout(w65_124));
	PE pe65_125(.x(x125),.w(w65_124),.acc(r65_124),.res(r65_125),.clk(clk),.wout(w65_125));
	PE pe65_126(.x(x126),.w(w65_125),.acc(r65_125),.res(r65_126),.clk(clk),.wout(w65_126));
	PE pe65_127(.x(x127),.w(w65_126),.acc(r65_126),.res(result65),.clk(clk),.wout(weight65));

	PE pe66_0(.x(x0),.w(w66),.acc(32'h0),.res(r66_0),.clk(clk),.wout(w66_0));
	PE pe66_1(.x(x1),.w(w66_0),.acc(r66_0),.res(r66_1),.clk(clk),.wout(w66_1));
	PE pe66_2(.x(x2),.w(w66_1),.acc(r66_1),.res(r66_2),.clk(clk),.wout(w66_2));
	PE pe66_3(.x(x3),.w(w66_2),.acc(r66_2),.res(r66_3),.clk(clk),.wout(w66_3));
	PE pe66_4(.x(x4),.w(w66_3),.acc(r66_3),.res(r66_4),.clk(clk),.wout(w66_4));
	PE pe66_5(.x(x5),.w(w66_4),.acc(r66_4),.res(r66_5),.clk(clk),.wout(w66_5));
	PE pe66_6(.x(x6),.w(w66_5),.acc(r66_5),.res(r66_6),.clk(clk),.wout(w66_6));
	PE pe66_7(.x(x7),.w(w66_6),.acc(r66_6),.res(r66_7),.clk(clk),.wout(w66_7));
	PE pe66_8(.x(x8),.w(w66_7),.acc(r66_7),.res(r66_8),.clk(clk),.wout(w66_8));
	PE pe66_9(.x(x9),.w(w66_8),.acc(r66_8),.res(r66_9),.clk(clk),.wout(w66_9));
	PE pe66_10(.x(x10),.w(w66_9),.acc(r66_9),.res(r66_10),.clk(clk),.wout(w66_10));
	PE pe66_11(.x(x11),.w(w66_10),.acc(r66_10),.res(r66_11),.clk(clk),.wout(w66_11));
	PE pe66_12(.x(x12),.w(w66_11),.acc(r66_11),.res(r66_12),.clk(clk),.wout(w66_12));
	PE pe66_13(.x(x13),.w(w66_12),.acc(r66_12),.res(r66_13),.clk(clk),.wout(w66_13));
	PE pe66_14(.x(x14),.w(w66_13),.acc(r66_13),.res(r66_14),.clk(clk),.wout(w66_14));
	PE pe66_15(.x(x15),.w(w66_14),.acc(r66_14),.res(r66_15),.clk(clk),.wout(w66_15));
	PE pe66_16(.x(x16),.w(w66_15),.acc(r66_15),.res(r66_16),.clk(clk),.wout(w66_16));
	PE pe66_17(.x(x17),.w(w66_16),.acc(r66_16),.res(r66_17),.clk(clk),.wout(w66_17));
	PE pe66_18(.x(x18),.w(w66_17),.acc(r66_17),.res(r66_18),.clk(clk),.wout(w66_18));
	PE pe66_19(.x(x19),.w(w66_18),.acc(r66_18),.res(r66_19),.clk(clk),.wout(w66_19));
	PE pe66_20(.x(x20),.w(w66_19),.acc(r66_19),.res(r66_20),.clk(clk),.wout(w66_20));
	PE pe66_21(.x(x21),.w(w66_20),.acc(r66_20),.res(r66_21),.clk(clk),.wout(w66_21));
	PE pe66_22(.x(x22),.w(w66_21),.acc(r66_21),.res(r66_22),.clk(clk),.wout(w66_22));
	PE pe66_23(.x(x23),.w(w66_22),.acc(r66_22),.res(r66_23),.clk(clk),.wout(w66_23));
	PE pe66_24(.x(x24),.w(w66_23),.acc(r66_23),.res(r66_24),.clk(clk),.wout(w66_24));
	PE pe66_25(.x(x25),.w(w66_24),.acc(r66_24),.res(r66_25),.clk(clk),.wout(w66_25));
	PE pe66_26(.x(x26),.w(w66_25),.acc(r66_25),.res(r66_26),.clk(clk),.wout(w66_26));
	PE pe66_27(.x(x27),.w(w66_26),.acc(r66_26),.res(r66_27),.clk(clk),.wout(w66_27));
	PE pe66_28(.x(x28),.w(w66_27),.acc(r66_27),.res(r66_28),.clk(clk),.wout(w66_28));
	PE pe66_29(.x(x29),.w(w66_28),.acc(r66_28),.res(r66_29),.clk(clk),.wout(w66_29));
	PE pe66_30(.x(x30),.w(w66_29),.acc(r66_29),.res(r66_30),.clk(clk),.wout(w66_30));
	PE pe66_31(.x(x31),.w(w66_30),.acc(r66_30),.res(r66_31),.clk(clk),.wout(w66_31));
	PE pe66_32(.x(x32),.w(w66_31),.acc(r66_31),.res(r66_32),.clk(clk),.wout(w66_32));
	PE pe66_33(.x(x33),.w(w66_32),.acc(r66_32),.res(r66_33),.clk(clk),.wout(w66_33));
	PE pe66_34(.x(x34),.w(w66_33),.acc(r66_33),.res(r66_34),.clk(clk),.wout(w66_34));
	PE pe66_35(.x(x35),.w(w66_34),.acc(r66_34),.res(r66_35),.clk(clk),.wout(w66_35));
	PE pe66_36(.x(x36),.w(w66_35),.acc(r66_35),.res(r66_36),.clk(clk),.wout(w66_36));
	PE pe66_37(.x(x37),.w(w66_36),.acc(r66_36),.res(r66_37),.clk(clk),.wout(w66_37));
	PE pe66_38(.x(x38),.w(w66_37),.acc(r66_37),.res(r66_38),.clk(clk),.wout(w66_38));
	PE pe66_39(.x(x39),.w(w66_38),.acc(r66_38),.res(r66_39),.clk(clk),.wout(w66_39));
	PE pe66_40(.x(x40),.w(w66_39),.acc(r66_39),.res(r66_40),.clk(clk),.wout(w66_40));
	PE pe66_41(.x(x41),.w(w66_40),.acc(r66_40),.res(r66_41),.clk(clk),.wout(w66_41));
	PE pe66_42(.x(x42),.w(w66_41),.acc(r66_41),.res(r66_42),.clk(clk),.wout(w66_42));
	PE pe66_43(.x(x43),.w(w66_42),.acc(r66_42),.res(r66_43),.clk(clk),.wout(w66_43));
	PE pe66_44(.x(x44),.w(w66_43),.acc(r66_43),.res(r66_44),.clk(clk),.wout(w66_44));
	PE pe66_45(.x(x45),.w(w66_44),.acc(r66_44),.res(r66_45),.clk(clk),.wout(w66_45));
	PE pe66_46(.x(x46),.w(w66_45),.acc(r66_45),.res(r66_46),.clk(clk),.wout(w66_46));
	PE pe66_47(.x(x47),.w(w66_46),.acc(r66_46),.res(r66_47),.clk(clk),.wout(w66_47));
	PE pe66_48(.x(x48),.w(w66_47),.acc(r66_47),.res(r66_48),.clk(clk),.wout(w66_48));
	PE pe66_49(.x(x49),.w(w66_48),.acc(r66_48),.res(r66_49),.clk(clk),.wout(w66_49));
	PE pe66_50(.x(x50),.w(w66_49),.acc(r66_49),.res(r66_50),.clk(clk),.wout(w66_50));
	PE pe66_51(.x(x51),.w(w66_50),.acc(r66_50),.res(r66_51),.clk(clk),.wout(w66_51));
	PE pe66_52(.x(x52),.w(w66_51),.acc(r66_51),.res(r66_52),.clk(clk),.wout(w66_52));
	PE pe66_53(.x(x53),.w(w66_52),.acc(r66_52),.res(r66_53),.clk(clk),.wout(w66_53));
	PE pe66_54(.x(x54),.w(w66_53),.acc(r66_53),.res(r66_54),.clk(clk),.wout(w66_54));
	PE pe66_55(.x(x55),.w(w66_54),.acc(r66_54),.res(r66_55),.clk(clk),.wout(w66_55));
	PE pe66_56(.x(x56),.w(w66_55),.acc(r66_55),.res(r66_56),.clk(clk),.wout(w66_56));
	PE pe66_57(.x(x57),.w(w66_56),.acc(r66_56),.res(r66_57),.clk(clk),.wout(w66_57));
	PE pe66_58(.x(x58),.w(w66_57),.acc(r66_57),.res(r66_58),.clk(clk),.wout(w66_58));
	PE pe66_59(.x(x59),.w(w66_58),.acc(r66_58),.res(r66_59),.clk(clk),.wout(w66_59));
	PE pe66_60(.x(x60),.w(w66_59),.acc(r66_59),.res(r66_60),.clk(clk),.wout(w66_60));
	PE pe66_61(.x(x61),.w(w66_60),.acc(r66_60),.res(r66_61),.clk(clk),.wout(w66_61));
	PE pe66_62(.x(x62),.w(w66_61),.acc(r66_61),.res(r66_62),.clk(clk),.wout(w66_62));
	PE pe66_63(.x(x63),.w(w66_62),.acc(r66_62),.res(r66_63),.clk(clk),.wout(w66_63));
	PE pe66_64(.x(x64),.w(w66_63),.acc(r66_63),.res(r66_64),.clk(clk),.wout(w66_64));
	PE pe66_65(.x(x65),.w(w66_64),.acc(r66_64),.res(r66_65),.clk(clk),.wout(w66_65));
	PE pe66_66(.x(x66),.w(w66_65),.acc(r66_65),.res(r66_66),.clk(clk),.wout(w66_66));
	PE pe66_67(.x(x67),.w(w66_66),.acc(r66_66),.res(r66_67),.clk(clk),.wout(w66_67));
	PE pe66_68(.x(x68),.w(w66_67),.acc(r66_67),.res(r66_68),.clk(clk),.wout(w66_68));
	PE pe66_69(.x(x69),.w(w66_68),.acc(r66_68),.res(r66_69),.clk(clk),.wout(w66_69));
	PE pe66_70(.x(x70),.w(w66_69),.acc(r66_69),.res(r66_70),.clk(clk),.wout(w66_70));
	PE pe66_71(.x(x71),.w(w66_70),.acc(r66_70),.res(r66_71),.clk(clk),.wout(w66_71));
	PE pe66_72(.x(x72),.w(w66_71),.acc(r66_71),.res(r66_72),.clk(clk),.wout(w66_72));
	PE pe66_73(.x(x73),.w(w66_72),.acc(r66_72),.res(r66_73),.clk(clk),.wout(w66_73));
	PE pe66_74(.x(x74),.w(w66_73),.acc(r66_73),.res(r66_74),.clk(clk),.wout(w66_74));
	PE pe66_75(.x(x75),.w(w66_74),.acc(r66_74),.res(r66_75),.clk(clk),.wout(w66_75));
	PE pe66_76(.x(x76),.w(w66_75),.acc(r66_75),.res(r66_76),.clk(clk),.wout(w66_76));
	PE pe66_77(.x(x77),.w(w66_76),.acc(r66_76),.res(r66_77),.clk(clk),.wout(w66_77));
	PE pe66_78(.x(x78),.w(w66_77),.acc(r66_77),.res(r66_78),.clk(clk),.wout(w66_78));
	PE pe66_79(.x(x79),.w(w66_78),.acc(r66_78),.res(r66_79),.clk(clk),.wout(w66_79));
	PE pe66_80(.x(x80),.w(w66_79),.acc(r66_79),.res(r66_80),.clk(clk),.wout(w66_80));
	PE pe66_81(.x(x81),.w(w66_80),.acc(r66_80),.res(r66_81),.clk(clk),.wout(w66_81));
	PE pe66_82(.x(x82),.w(w66_81),.acc(r66_81),.res(r66_82),.clk(clk),.wout(w66_82));
	PE pe66_83(.x(x83),.w(w66_82),.acc(r66_82),.res(r66_83),.clk(clk),.wout(w66_83));
	PE pe66_84(.x(x84),.w(w66_83),.acc(r66_83),.res(r66_84),.clk(clk),.wout(w66_84));
	PE pe66_85(.x(x85),.w(w66_84),.acc(r66_84),.res(r66_85),.clk(clk),.wout(w66_85));
	PE pe66_86(.x(x86),.w(w66_85),.acc(r66_85),.res(r66_86),.clk(clk),.wout(w66_86));
	PE pe66_87(.x(x87),.w(w66_86),.acc(r66_86),.res(r66_87),.clk(clk),.wout(w66_87));
	PE pe66_88(.x(x88),.w(w66_87),.acc(r66_87),.res(r66_88),.clk(clk),.wout(w66_88));
	PE pe66_89(.x(x89),.w(w66_88),.acc(r66_88),.res(r66_89),.clk(clk),.wout(w66_89));
	PE pe66_90(.x(x90),.w(w66_89),.acc(r66_89),.res(r66_90),.clk(clk),.wout(w66_90));
	PE pe66_91(.x(x91),.w(w66_90),.acc(r66_90),.res(r66_91),.clk(clk),.wout(w66_91));
	PE pe66_92(.x(x92),.w(w66_91),.acc(r66_91),.res(r66_92),.clk(clk),.wout(w66_92));
	PE pe66_93(.x(x93),.w(w66_92),.acc(r66_92),.res(r66_93),.clk(clk),.wout(w66_93));
	PE pe66_94(.x(x94),.w(w66_93),.acc(r66_93),.res(r66_94),.clk(clk),.wout(w66_94));
	PE pe66_95(.x(x95),.w(w66_94),.acc(r66_94),.res(r66_95),.clk(clk),.wout(w66_95));
	PE pe66_96(.x(x96),.w(w66_95),.acc(r66_95),.res(r66_96),.clk(clk),.wout(w66_96));
	PE pe66_97(.x(x97),.w(w66_96),.acc(r66_96),.res(r66_97),.clk(clk),.wout(w66_97));
	PE pe66_98(.x(x98),.w(w66_97),.acc(r66_97),.res(r66_98),.clk(clk),.wout(w66_98));
	PE pe66_99(.x(x99),.w(w66_98),.acc(r66_98),.res(r66_99),.clk(clk),.wout(w66_99));
	PE pe66_100(.x(x100),.w(w66_99),.acc(r66_99),.res(r66_100),.clk(clk),.wout(w66_100));
	PE pe66_101(.x(x101),.w(w66_100),.acc(r66_100),.res(r66_101),.clk(clk),.wout(w66_101));
	PE pe66_102(.x(x102),.w(w66_101),.acc(r66_101),.res(r66_102),.clk(clk),.wout(w66_102));
	PE pe66_103(.x(x103),.w(w66_102),.acc(r66_102),.res(r66_103),.clk(clk),.wout(w66_103));
	PE pe66_104(.x(x104),.w(w66_103),.acc(r66_103),.res(r66_104),.clk(clk),.wout(w66_104));
	PE pe66_105(.x(x105),.w(w66_104),.acc(r66_104),.res(r66_105),.clk(clk),.wout(w66_105));
	PE pe66_106(.x(x106),.w(w66_105),.acc(r66_105),.res(r66_106),.clk(clk),.wout(w66_106));
	PE pe66_107(.x(x107),.w(w66_106),.acc(r66_106),.res(r66_107),.clk(clk),.wout(w66_107));
	PE pe66_108(.x(x108),.w(w66_107),.acc(r66_107),.res(r66_108),.clk(clk),.wout(w66_108));
	PE pe66_109(.x(x109),.w(w66_108),.acc(r66_108),.res(r66_109),.clk(clk),.wout(w66_109));
	PE pe66_110(.x(x110),.w(w66_109),.acc(r66_109),.res(r66_110),.clk(clk),.wout(w66_110));
	PE pe66_111(.x(x111),.w(w66_110),.acc(r66_110),.res(r66_111),.clk(clk),.wout(w66_111));
	PE pe66_112(.x(x112),.w(w66_111),.acc(r66_111),.res(r66_112),.clk(clk),.wout(w66_112));
	PE pe66_113(.x(x113),.w(w66_112),.acc(r66_112),.res(r66_113),.clk(clk),.wout(w66_113));
	PE pe66_114(.x(x114),.w(w66_113),.acc(r66_113),.res(r66_114),.clk(clk),.wout(w66_114));
	PE pe66_115(.x(x115),.w(w66_114),.acc(r66_114),.res(r66_115),.clk(clk),.wout(w66_115));
	PE pe66_116(.x(x116),.w(w66_115),.acc(r66_115),.res(r66_116),.clk(clk),.wout(w66_116));
	PE pe66_117(.x(x117),.w(w66_116),.acc(r66_116),.res(r66_117),.clk(clk),.wout(w66_117));
	PE pe66_118(.x(x118),.w(w66_117),.acc(r66_117),.res(r66_118),.clk(clk),.wout(w66_118));
	PE pe66_119(.x(x119),.w(w66_118),.acc(r66_118),.res(r66_119),.clk(clk),.wout(w66_119));
	PE pe66_120(.x(x120),.w(w66_119),.acc(r66_119),.res(r66_120),.clk(clk),.wout(w66_120));
	PE pe66_121(.x(x121),.w(w66_120),.acc(r66_120),.res(r66_121),.clk(clk),.wout(w66_121));
	PE pe66_122(.x(x122),.w(w66_121),.acc(r66_121),.res(r66_122),.clk(clk),.wout(w66_122));
	PE pe66_123(.x(x123),.w(w66_122),.acc(r66_122),.res(r66_123),.clk(clk),.wout(w66_123));
	PE pe66_124(.x(x124),.w(w66_123),.acc(r66_123),.res(r66_124),.clk(clk),.wout(w66_124));
	PE pe66_125(.x(x125),.w(w66_124),.acc(r66_124),.res(r66_125),.clk(clk),.wout(w66_125));
	PE pe66_126(.x(x126),.w(w66_125),.acc(r66_125),.res(r66_126),.clk(clk),.wout(w66_126));
	PE pe66_127(.x(x127),.w(w66_126),.acc(r66_126),.res(result66),.clk(clk),.wout(weight66));

	PE pe67_0(.x(x0),.w(w67),.acc(32'h0),.res(r67_0),.clk(clk),.wout(w67_0));
	PE pe67_1(.x(x1),.w(w67_0),.acc(r67_0),.res(r67_1),.clk(clk),.wout(w67_1));
	PE pe67_2(.x(x2),.w(w67_1),.acc(r67_1),.res(r67_2),.clk(clk),.wout(w67_2));
	PE pe67_3(.x(x3),.w(w67_2),.acc(r67_2),.res(r67_3),.clk(clk),.wout(w67_3));
	PE pe67_4(.x(x4),.w(w67_3),.acc(r67_3),.res(r67_4),.clk(clk),.wout(w67_4));
	PE pe67_5(.x(x5),.w(w67_4),.acc(r67_4),.res(r67_5),.clk(clk),.wout(w67_5));
	PE pe67_6(.x(x6),.w(w67_5),.acc(r67_5),.res(r67_6),.clk(clk),.wout(w67_6));
	PE pe67_7(.x(x7),.w(w67_6),.acc(r67_6),.res(r67_7),.clk(clk),.wout(w67_7));
	PE pe67_8(.x(x8),.w(w67_7),.acc(r67_7),.res(r67_8),.clk(clk),.wout(w67_8));
	PE pe67_9(.x(x9),.w(w67_8),.acc(r67_8),.res(r67_9),.clk(clk),.wout(w67_9));
	PE pe67_10(.x(x10),.w(w67_9),.acc(r67_9),.res(r67_10),.clk(clk),.wout(w67_10));
	PE pe67_11(.x(x11),.w(w67_10),.acc(r67_10),.res(r67_11),.clk(clk),.wout(w67_11));
	PE pe67_12(.x(x12),.w(w67_11),.acc(r67_11),.res(r67_12),.clk(clk),.wout(w67_12));
	PE pe67_13(.x(x13),.w(w67_12),.acc(r67_12),.res(r67_13),.clk(clk),.wout(w67_13));
	PE pe67_14(.x(x14),.w(w67_13),.acc(r67_13),.res(r67_14),.clk(clk),.wout(w67_14));
	PE pe67_15(.x(x15),.w(w67_14),.acc(r67_14),.res(r67_15),.clk(clk),.wout(w67_15));
	PE pe67_16(.x(x16),.w(w67_15),.acc(r67_15),.res(r67_16),.clk(clk),.wout(w67_16));
	PE pe67_17(.x(x17),.w(w67_16),.acc(r67_16),.res(r67_17),.clk(clk),.wout(w67_17));
	PE pe67_18(.x(x18),.w(w67_17),.acc(r67_17),.res(r67_18),.clk(clk),.wout(w67_18));
	PE pe67_19(.x(x19),.w(w67_18),.acc(r67_18),.res(r67_19),.clk(clk),.wout(w67_19));
	PE pe67_20(.x(x20),.w(w67_19),.acc(r67_19),.res(r67_20),.clk(clk),.wout(w67_20));
	PE pe67_21(.x(x21),.w(w67_20),.acc(r67_20),.res(r67_21),.clk(clk),.wout(w67_21));
	PE pe67_22(.x(x22),.w(w67_21),.acc(r67_21),.res(r67_22),.clk(clk),.wout(w67_22));
	PE pe67_23(.x(x23),.w(w67_22),.acc(r67_22),.res(r67_23),.clk(clk),.wout(w67_23));
	PE pe67_24(.x(x24),.w(w67_23),.acc(r67_23),.res(r67_24),.clk(clk),.wout(w67_24));
	PE pe67_25(.x(x25),.w(w67_24),.acc(r67_24),.res(r67_25),.clk(clk),.wout(w67_25));
	PE pe67_26(.x(x26),.w(w67_25),.acc(r67_25),.res(r67_26),.clk(clk),.wout(w67_26));
	PE pe67_27(.x(x27),.w(w67_26),.acc(r67_26),.res(r67_27),.clk(clk),.wout(w67_27));
	PE pe67_28(.x(x28),.w(w67_27),.acc(r67_27),.res(r67_28),.clk(clk),.wout(w67_28));
	PE pe67_29(.x(x29),.w(w67_28),.acc(r67_28),.res(r67_29),.clk(clk),.wout(w67_29));
	PE pe67_30(.x(x30),.w(w67_29),.acc(r67_29),.res(r67_30),.clk(clk),.wout(w67_30));
	PE pe67_31(.x(x31),.w(w67_30),.acc(r67_30),.res(r67_31),.clk(clk),.wout(w67_31));
	PE pe67_32(.x(x32),.w(w67_31),.acc(r67_31),.res(r67_32),.clk(clk),.wout(w67_32));
	PE pe67_33(.x(x33),.w(w67_32),.acc(r67_32),.res(r67_33),.clk(clk),.wout(w67_33));
	PE pe67_34(.x(x34),.w(w67_33),.acc(r67_33),.res(r67_34),.clk(clk),.wout(w67_34));
	PE pe67_35(.x(x35),.w(w67_34),.acc(r67_34),.res(r67_35),.clk(clk),.wout(w67_35));
	PE pe67_36(.x(x36),.w(w67_35),.acc(r67_35),.res(r67_36),.clk(clk),.wout(w67_36));
	PE pe67_37(.x(x37),.w(w67_36),.acc(r67_36),.res(r67_37),.clk(clk),.wout(w67_37));
	PE pe67_38(.x(x38),.w(w67_37),.acc(r67_37),.res(r67_38),.clk(clk),.wout(w67_38));
	PE pe67_39(.x(x39),.w(w67_38),.acc(r67_38),.res(r67_39),.clk(clk),.wout(w67_39));
	PE pe67_40(.x(x40),.w(w67_39),.acc(r67_39),.res(r67_40),.clk(clk),.wout(w67_40));
	PE pe67_41(.x(x41),.w(w67_40),.acc(r67_40),.res(r67_41),.clk(clk),.wout(w67_41));
	PE pe67_42(.x(x42),.w(w67_41),.acc(r67_41),.res(r67_42),.clk(clk),.wout(w67_42));
	PE pe67_43(.x(x43),.w(w67_42),.acc(r67_42),.res(r67_43),.clk(clk),.wout(w67_43));
	PE pe67_44(.x(x44),.w(w67_43),.acc(r67_43),.res(r67_44),.clk(clk),.wout(w67_44));
	PE pe67_45(.x(x45),.w(w67_44),.acc(r67_44),.res(r67_45),.clk(clk),.wout(w67_45));
	PE pe67_46(.x(x46),.w(w67_45),.acc(r67_45),.res(r67_46),.clk(clk),.wout(w67_46));
	PE pe67_47(.x(x47),.w(w67_46),.acc(r67_46),.res(r67_47),.clk(clk),.wout(w67_47));
	PE pe67_48(.x(x48),.w(w67_47),.acc(r67_47),.res(r67_48),.clk(clk),.wout(w67_48));
	PE pe67_49(.x(x49),.w(w67_48),.acc(r67_48),.res(r67_49),.clk(clk),.wout(w67_49));
	PE pe67_50(.x(x50),.w(w67_49),.acc(r67_49),.res(r67_50),.clk(clk),.wout(w67_50));
	PE pe67_51(.x(x51),.w(w67_50),.acc(r67_50),.res(r67_51),.clk(clk),.wout(w67_51));
	PE pe67_52(.x(x52),.w(w67_51),.acc(r67_51),.res(r67_52),.clk(clk),.wout(w67_52));
	PE pe67_53(.x(x53),.w(w67_52),.acc(r67_52),.res(r67_53),.clk(clk),.wout(w67_53));
	PE pe67_54(.x(x54),.w(w67_53),.acc(r67_53),.res(r67_54),.clk(clk),.wout(w67_54));
	PE pe67_55(.x(x55),.w(w67_54),.acc(r67_54),.res(r67_55),.clk(clk),.wout(w67_55));
	PE pe67_56(.x(x56),.w(w67_55),.acc(r67_55),.res(r67_56),.clk(clk),.wout(w67_56));
	PE pe67_57(.x(x57),.w(w67_56),.acc(r67_56),.res(r67_57),.clk(clk),.wout(w67_57));
	PE pe67_58(.x(x58),.w(w67_57),.acc(r67_57),.res(r67_58),.clk(clk),.wout(w67_58));
	PE pe67_59(.x(x59),.w(w67_58),.acc(r67_58),.res(r67_59),.clk(clk),.wout(w67_59));
	PE pe67_60(.x(x60),.w(w67_59),.acc(r67_59),.res(r67_60),.clk(clk),.wout(w67_60));
	PE pe67_61(.x(x61),.w(w67_60),.acc(r67_60),.res(r67_61),.clk(clk),.wout(w67_61));
	PE pe67_62(.x(x62),.w(w67_61),.acc(r67_61),.res(r67_62),.clk(clk),.wout(w67_62));
	PE pe67_63(.x(x63),.w(w67_62),.acc(r67_62),.res(r67_63),.clk(clk),.wout(w67_63));
	PE pe67_64(.x(x64),.w(w67_63),.acc(r67_63),.res(r67_64),.clk(clk),.wout(w67_64));
	PE pe67_65(.x(x65),.w(w67_64),.acc(r67_64),.res(r67_65),.clk(clk),.wout(w67_65));
	PE pe67_66(.x(x66),.w(w67_65),.acc(r67_65),.res(r67_66),.clk(clk),.wout(w67_66));
	PE pe67_67(.x(x67),.w(w67_66),.acc(r67_66),.res(r67_67),.clk(clk),.wout(w67_67));
	PE pe67_68(.x(x68),.w(w67_67),.acc(r67_67),.res(r67_68),.clk(clk),.wout(w67_68));
	PE pe67_69(.x(x69),.w(w67_68),.acc(r67_68),.res(r67_69),.clk(clk),.wout(w67_69));
	PE pe67_70(.x(x70),.w(w67_69),.acc(r67_69),.res(r67_70),.clk(clk),.wout(w67_70));
	PE pe67_71(.x(x71),.w(w67_70),.acc(r67_70),.res(r67_71),.clk(clk),.wout(w67_71));
	PE pe67_72(.x(x72),.w(w67_71),.acc(r67_71),.res(r67_72),.clk(clk),.wout(w67_72));
	PE pe67_73(.x(x73),.w(w67_72),.acc(r67_72),.res(r67_73),.clk(clk),.wout(w67_73));
	PE pe67_74(.x(x74),.w(w67_73),.acc(r67_73),.res(r67_74),.clk(clk),.wout(w67_74));
	PE pe67_75(.x(x75),.w(w67_74),.acc(r67_74),.res(r67_75),.clk(clk),.wout(w67_75));
	PE pe67_76(.x(x76),.w(w67_75),.acc(r67_75),.res(r67_76),.clk(clk),.wout(w67_76));
	PE pe67_77(.x(x77),.w(w67_76),.acc(r67_76),.res(r67_77),.clk(clk),.wout(w67_77));
	PE pe67_78(.x(x78),.w(w67_77),.acc(r67_77),.res(r67_78),.clk(clk),.wout(w67_78));
	PE pe67_79(.x(x79),.w(w67_78),.acc(r67_78),.res(r67_79),.clk(clk),.wout(w67_79));
	PE pe67_80(.x(x80),.w(w67_79),.acc(r67_79),.res(r67_80),.clk(clk),.wout(w67_80));
	PE pe67_81(.x(x81),.w(w67_80),.acc(r67_80),.res(r67_81),.clk(clk),.wout(w67_81));
	PE pe67_82(.x(x82),.w(w67_81),.acc(r67_81),.res(r67_82),.clk(clk),.wout(w67_82));
	PE pe67_83(.x(x83),.w(w67_82),.acc(r67_82),.res(r67_83),.clk(clk),.wout(w67_83));
	PE pe67_84(.x(x84),.w(w67_83),.acc(r67_83),.res(r67_84),.clk(clk),.wout(w67_84));
	PE pe67_85(.x(x85),.w(w67_84),.acc(r67_84),.res(r67_85),.clk(clk),.wout(w67_85));
	PE pe67_86(.x(x86),.w(w67_85),.acc(r67_85),.res(r67_86),.clk(clk),.wout(w67_86));
	PE pe67_87(.x(x87),.w(w67_86),.acc(r67_86),.res(r67_87),.clk(clk),.wout(w67_87));
	PE pe67_88(.x(x88),.w(w67_87),.acc(r67_87),.res(r67_88),.clk(clk),.wout(w67_88));
	PE pe67_89(.x(x89),.w(w67_88),.acc(r67_88),.res(r67_89),.clk(clk),.wout(w67_89));
	PE pe67_90(.x(x90),.w(w67_89),.acc(r67_89),.res(r67_90),.clk(clk),.wout(w67_90));
	PE pe67_91(.x(x91),.w(w67_90),.acc(r67_90),.res(r67_91),.clk(clk),.wout(w67_91));
	PE pe67_92(.x(x92),.w(w67_91),.acc(r67_91),.res(r67_92),.clk(clk),.wout(w67_92));
	PE pe67_93(.x(x93),.w(w67_92),.acc(r67_92),.res(r67_93),.clk(clk),.wout(w67_93));
	PE pe67_94(.x(x94),.w(w67_93),.acc(r67_93),.res(r67_94),.clk(clk),.wout(w67_94));
	PE pe67_95(.x(x95),.w(w67_94),.acc(r67_94),.res(r67_95),.clk(clk),.wout(w67_95));
	PE pe67_96(.x(x96),.w(w67_95),.acc(r67_95),.res(r67_96),.clk(clk),.wout(w67_96));
	PE pe67_97(.x(x97),.w(w67_96),.acc(r67_96),.res(r67_97),.clk(clk),.wout(w67_97));
	PE pe67_98(.x(x98),.w(w67_97),.acc(r67_97),.res(r67_98),.clk(clk),.wout(w67_98));
	PE pe67_99(.x(x99),.w(w67_98),.acc(r67_98),.res(r67_99),.clk(clk),.wout(w67_99));
	PE pe67_100(.x(x100),.w(w67_99),.acc(r67_99),.res(r67_100),.clk(clk),.wout(w67_100));
	PE pe67_101(.x(x101),.w(w67_100),.acc(r67_100),.res(r67_101),.clk(clk),.wout(w67_101));
	PE pe67_102(.x(x102),.w(w67_101),.acc(r67_101),.res(r67_102),.clk(clk),.wout(w67_102));
	PE pe67_103(.x(x103),.w(w67_102),.acc(r67_102),.res(r67_103),.clk(clk),.wout(w67_103));
	PE pe67_104(.x(x104),.w(w67_103),.acc(r67_103),.res(r67_104),.clk(clk),.wout(w67_104));
	PE pe67_105(.x(x105),.w(w67_104),.acc(r67_104),.res(r67_105),.clk(clk),.wout(w67_105));
	PE pe67_106(.x(x106),.w(w67_105),.acc(r67_105),.res(r67_106),.clk(clk),.wout(w67_106));
	PE pe67_107(.x(x107),.w(w67_106),.acc(r67_106),.res(r67_107),.clk(clk),.wout(w67_107));
	PE pe67_108(.x(x108),.w(w67_107),.acc(r67_107),.res(r67_108),.clk(clk),.wout(w67_108));
	PE pe67_109(.x(x109),.w(w67_108),.acc(r67_108),.res(r67_109),.clk(clk),.wout(w67_109));
	PE pe67_110(.x(x110),.w(w67_109),.acc(r67_109),.res(r67_110),.clk(clk),.wout(w67_110));
	PE pe67_111(.x(x111),.w(w67_110),.acc(r67_110),.res(r67_111),.clk(clk),.wout(w67_111));
	PE pe67_112(.x(x112),.w(w67_111),.acc(r67_111),.res(r67_112),.clk(clk),.wout(w67_112));
	PE pe67_113(.x(x113),.w(w67_112),.acc(r67_112),.res(r67_113),.clk(clk),.wout(w67_113));
	PE pe67_114(.x(x114),.w(w67_113),.acc(r67_113),.res(r67_114),.clk(clk),.wout(w67_114));
	PE pe67_115(.x(x115),.w(w67_114),.acc(r67_114),.res(r67_115),.clk(clk),.wout(w67_115));
	PE pe67_116(.x(x116),.w(w67_115),.acc(r67_115),.res(r67_116),.clk(clk),.wout(w67_116));
	PE pe67_117(.x(x117),.w(w67_116),.acc(r67_116),.res(r67_117),.clk(clk),.wout(w67_117));
	PE pe67_118(.x(x118),.w(w67_117),.acc(r67_117),.res(r67_118),.clk(clk),.wout(w67_118));
	PE pe67_119(.x(x119),.w(w67_118),.acc(r67_118),.res(r67_119),.clk(clk),.wout(w67_119));
	PE pe67_120(.x(x120),.w(w67_119),.acc(r67_119),.res(r67_120),.clk(clk),.wout(w67_120));
	PE pe67_121(.x(x121),.w(w67_120),.acc(r67_120),.res(r67_121),.clk(clk),.wout(w67_121));
	PE pe67_122(.x(x122),.w(w67_121),.acc(r67_121),.res(r67_122),.clk(clk),.wout(w67_122));
	PE pe67_123(.x(x123),.w(w67_122),.acc(r67_122),.res(r67_123),.clk(clk),.wout(w67_123));
	PE pe67_124(.x(x124),.w(w67_123),.acc(r67_123),.res(r67_124),.clk(clk),.wout(w67_124));
	PE pe67_125(.x(x125),.w(w67_124),.acc(r67_124),.res(r67_125),.clk(clk),.wout(w67_125));
	PE pe67_126(.x(x126),.w(w67_125),.acc(r67_125),.res(r67_126),.clk(clk),.wout(w67_126));
	PE pe67_127(.x(x127),.w(w67_126),.acc(r67_126),.res(result67),.clk(clk),.wout(weight67));

	PE pe68_0(.x(x0),.w(w68),.acc(32'h0),.res(r68_0),.clk(clk),.wout(w68_0));
	PE pe68_1(.x(x1),.w(w68_0),.acc(r68_0),.res(r68_1),.clk(clk),.wout(w68_1));
	PE pe68_2(.x(x2),.w(w68_1),.acc(r68_1),.res(r68_2),.clk(clk),.wout(w68_2));
	PE pe68_3(.x(x3),.w(w68_2),.acc(r68_2),.res(r68_3),.clk(clk),.wout(w68_3));
	PE pe68_4(.x(x4),.w(w68_3),.acc(r68_3),.res(r68_4),.clk(clk),.wout(w68_4));
	PE pe68_5(.x(x5),.w(w68_4),.acc(r68_4),.res(r68_5),.clk(clk),.wout(w68_5));
	PE pe68_6(.x(x6),.w(w68_5),.acc(r68_5),.res(r68_6),.clk(clk),.wout(w68_6));
	PE pe68_7(.x(x7),.w(w68_6),.acc(r68_6),.res(r68_7),.clk(clk),.wout(w68_7));
	PE pe68_8(.x(x8),.w(w68_7),.acc(r68_7),.res(r68_8),.clk(clk),.wout(w68_8));
	PE pe68_9(.x(x9),.w(w68_8),.acc(r68_8),.res(r68_9),.clk(clk),.wout(w68_9));
	PE pe68_10(.x(x10),.w(w68_9),.acc(r68_9),.res(r68_10),.clk(clk),.wout(w68_10));
	PE pe68_11(.x(x11),.w(w68_10),.acc(r68_10),.res(r68_11),.clk(clk),.wout(w68_11));
	PE pe68_12(.x(x12),.w(w68_11),.acc(r68_11),.res(r68_12),.clk(clk),.wout(w68_12));
	PE pe68_13(.x(x13),.w(w68_12),.acc(r68_12),.res(r68_13),.clk(clk),.wout(w68_13));
	PE pe68_14(.x(x14),.w(w68_13),.acc(r68_13),.res(r68_14),.clk(clk),.wout(w68_14));
	PE pe68_15(.x(x15),.w(w68_14),.acc(r68_14),.res(r68_15),.clk(clk),.wout(w68_15));
	PE pe68_16(.x(x16),.w(w68_15),.acc(r68_15),.res(r68_16),.clk(clk),.wout(w68_16));
	PE pe68_17(.x(x17),.w(w68_16),.acc(r68_16),.res(r68_17),.clk(clk),.wout(w68_17));
	PE pe68_18(.x(x18),.w(w68_17),.acc(r68_17),.res(r68_18),.clk(clk),.wout(w68_18));
	PE pe68_19(.x(x19),.w(w68_18),.acc(r68_18),.res(r68_19),.clk(clk),.wout(w68_19));
	PE pe68_20(.x(x20),.w(w68_19),.acc(r68_19),.res(r68_20),.clk(clk),.wout(w68_20));
	PE pe68_21(.x(x21),.w(w68_20),.acc(r68_20),.res(r68_21),.clk(clk),.wout(w68_21));
	PE pe68_22(.x(x22),.w(w68_21),.acc(r68_21),.res(r68_22),.clk(clk),.wout(w68_22));
	PE pe68_23(.x(x23),.w(w68_22),.acc(r68_22),.res(r68_23),.clk(clk),.wout(w68_23));
	PE pe68_24(.x(x24),.w(w68_23),.acc(r68_23),.res(r68_24),.clk(clk),.wout(w68_24));
	PE pe68_25(.x(x25),.w(w68_24),.acc(r68_24),.res(r68_25),.clk(clk),.wout(w68_25));
	PE pe68_26(.x(x26),.w(w68_25),.acc(r68_25),.res(r68_26),.clk(clk),.wout(w68_26));
	PE pe68_27(.x(x27),.w(w68_26),.acc(r68_26),.res(r68_27),.clk(clk),.wout(w68_27));
	PE pe68_28(.x(x28),.w(w68_27),.acc(r68_27),.res(r68_28),.clk(clk),.wout(w68_28));
	PE pe68_29(.x(x29),.w(w68_28),.acc(r68_28),.res(r68_29),.clk(clk),.wout(w68_29));
	PE pe68_30(.x(x30),.w(w68_29),.acc(r68_29),.res(r68_30),.clk(clk),.wout(w68_30));
	PE pe68_31(.x(x31),.w(w68_30),.acc(r68_30),.res(r68_31),.clk(clk),.wout(w68_31));
	PE pe68_32(.x(x32),.w(w68_31),.acc(r68_31),.res(r68_32),.clk(clk),.wout(w68_32));
	PE pe68_33(.x(x33),.w(w68_32),.acc(r68_32),.res(r68_33),.clk(clk),.wout(w68_33));
	PE pe68_34(.x(x34),.w(w68_33),.acc(r68_33),.res(r68_34),.clk(clk),.wout(w68_34));
	PE pe68_35(.x(x35),.w(w68_34),.acc(r68_34),.res(r68_35),.clk(clk),.wout(w68_35));
	PE pe68_36(.x(x36),.w(w68_35),.acc(r68_35),.res(r68_36),.clk(clk),.wout(w68_36));
	PE pe68_37(.x(x37),.w(w68_36),.acc(r68_36),.res(r68_37),.clk(clk),.wout(w68_37));
	PE pe68_38(.x(x38),.w(w68_37),.acc(r68_37),.res(r68_38),.clk(clk),.wout(w68_38));
	PE pe68_39(.x(x39),.w(w68_38),.acc(r68_38),.res(r68_39),.clk(clk),.wout(w68_39));
	PE pe68_40(.x(x40),.w(w68_39),.acc(r68_39),.res(r68_40),.clk(clk),.wout(w68_40));
	PE pe68_41(.x(x41),.w(w68_40),.acc(r68_40),.res(r68_41),.clk(clk),.wout(w68_41));
	PE pe68_42(.x(x42),.w(w68_41),.acc(r68_41),.res(r68_42),.clk(clk),.wout(w68_42));
	PE pe68_43(.x(x43),.w(w68_42),.acc(r68_42),.res(r68_43),.clk(clk),.wout(w68_43));
	PE pe68_44(.x(x44),.w(w68_43),.acc(r68_43),.res(r68_44),.clk(clk),.wout(w68_44));
	PE pe68_45(.x(x45),.w(w68_44),.acc(r68_44),.res(r68_45),.clk(clk),.wout(w68_45));
	PE pe68_46(.x(x46),.w(w68_45),.acc(r68_45),.res(r68_46),.clk(clk),.wout(w68_46));
	PE pe68_47(.x(x47),.w(w68_46),.acc(r68_46),.res(r68_47),.clk(clk),.wout(w68_47));
	PE pe68_48(.x(x48),.w(w68_47),.acc(r68_47),.res(r68_48),.clk(clk),.wout(w68_48));
	PE pe68_49(.x(x49),.w(w68_48),.acc(r68_48),.res(r68_49),.clk(clk),.wout(w68_49));
	PE pe68_50(.x(x50),.w(w68_49),.acc(r68_49),.res(r68_50),.clk(clk),.wout(w68_50));
	PE pe68_51(.x(x51),.w(w68_50),.acc(r68_50),.res(r68_51),.clk(clk),.wout(w68_51));
	PE pe68_52(.x(x52),.w(w68_51),.acc(r68_51),.res(r68_52),.clk(clk),.wout(w68_52));
	PE pe68_53(.x(x53),.w(w68_52),.acc(r68_52),.res(r68_53),.clk(clk),.wout(w68_53));
	PE pe68_54(.x(x54),.w(w68_53),.acc(r68_53),.res(r68_54),.clk(clk),.wout(w68_54));
	PE pe68_55(.x(x55),.w(w68_54),.acc(r68_54),.res(r68_55),.clk(clk),.wout(w68_55));
	PE pe68_56(.x(x56),.w(w68_55),.acc(r68_55),.res(r68_56),.clk(clk),.wout(w68_56));
	PE pe68_57(.x(x57),.w(w68_56),.acc(r68_56),.res(r68_57),.clk(clk),.wout(w68_57));
	PE pe68_58(.x(x58),.w(w68_57),.acc(r68_57),.res(r68_58),.clk(clk),.wout(w68_58));
	PE pe68_59(.x(x59),.w(w68_58),.acc(r68_58),.res(r68_59),.clk(clk),.wout(w68_59));
	PE pe68_60(.x(x60),.w(w68_59),.acc(r68_59),.res(r68_60),.clk(clk),.wout(w68_60));
	PE pe68_61(.x(x61),.w(w68_60),.acc(r68_60),.res(r68_61),.clk(clk),.wout(w68_61));
	PE pe68_62(.x(x62),.w(w68_61),.acc(r68_61),.res(r68_62),.clk(clk),.wout(w68_62));
	PE pe68_63(.x(x63),.w(w68_62),.acc(r68_62),.res(r68_63),.clk(clk),.wout(w68_63));
	PE pe68_64(.x(x64),.w(w68_63),.acc(r68_63),.res(r68_64),.clk(clk),.wout(w68_64));
	PE pe68_65(.x(x65),.w(w68_64),.acc(r68_64),.res(r68_65),.clk(clk),.wout(w68_65));
	PE pe68_66(.x(x66),.w(w68_65),.acc(r68_65),.res(r68_66),.clk(clk),.wout(w68_66));
	PE pe68_67(.x(x67),.w(w68_66),.acc(r68_66),.res(r68_67),.clk(clk),.wout(w68_67));
	PE pe68_68(.x(x68),.w(w68_67),.acc(r68_67),.res(r68_68),.clk(clk),.wout(w68_68));
	PE pe68_69(.x(x69),.w(w68_68),.acc(r68_68),.res(r68_69),.clk(clk),.wout(w68_69));
	PE pe68_70(.x(x70),.w(w68_69),.acc(r68_69),.res(r68_70),.clk(clk),.wout(w68_70));
	PE pe68_71(.x(x71),.w(w68_70),.acc(r68_70),.res(r68_71),.clk(clk),.wout(w68_71));
	PE pe68_72(.x(x72),.w(w68_71),.acc(r68_71),.res(r68_72),.clk(clk),.wout(w68_72));
	PE pe68_73(.x(x73),.w(w68_72),.acc(r68_72),.res(r68_73),.clk(clk),.wout(w68_73));
	PE pe68_74(.x(x74),.w(w68_73),.acc(r68_73),.res(r68_74),.clk(clk),.wout(w68_74));
	PE pe68_75(.x(x75),.w(w68_74),.acc(r68_74),.res(r68_75),.clk(clk),.wout(w68_75));
	PE pe68_76(.x(x76),.w(w68_75),.acc(r68_75),.res(r68_76),.clk(clk),.wout(w68_76));
	PE pe68_77(.x(x77),.w(w68_76),.acc(r68_76),.res(r68_77),.clk(clk),.wout(w68_77));
	PE pe68_78(.x(x78),.w(w68_77),.acc(r68_77),.res(r68_78),.clk(clk),.wout(w68_78));
	PE pe68_79(.x(x79),.w(w68_78),.acc(r68_78),.res(r68_79),.clk(clk),.wout(w68_79));
	PE pe68_80(.x(x80),.w(w68_79),.acc(r68_79),.res(r68_80),.clk(clk),.wout(w68_80));
	PE pe68_81(.x(x81),.w(w68_80),.acc(r68_80),.res(r68_81),.clk(clk),.wout(w68_81));
	PE pe68_82(.x(x82),.w(w68_81),.acc(r68_81),.res(r68_82),.clk(clk),.wout(w68_82));
	PE pe68_83(.x(x83),.w(w68_82),.acc(r68_82),.res(r68_83),.clk(clk),.wout(w68_83));
	PE pe68_84(.x(x84),.w(w68_83),.acc(r68_83),.res(r68_84),.clk(clk),.wout(w68_84));
	PE pe68_85(.x(x85),.w(w68_84),.acc(r68_84),.res(r68_85),.clk(clk),.wout(w68_85));
	PE pe68_86(.x(x86),.w(w68_85),.acc(r68_85),.res(r68_86),.clk(clk),.wout(w68_86));
	PE pe68_87(.x(x87),.w(w68_86),.acc(r68_86),.res(r68_87),.clk(clk),.wout(w68_87));
	PE pe68_88(.x(x88),.w(w68_87),.acc(r68_87),.res(r68_88),.clk(clk),.wout(w68_88));
	PE pe68_89(.x(x89),.w(w68_88),.acc(r68_88),.res(r68_89),.clk(clk),.wout(w68_89));
	PE pe68_90(.x(x90),.w(w68_89),.acc(r68_89),.res(r68_90),.clk(clk),.wout(w68_90));
	PE pe68_91(.x(x91),.w(w68_90),.acc(r68_90),.res(r68_91),.clk(clk),.wout(w68_91));
	PE pe68_92(.x(x92),.w(w68_91),.acc(r68_91),.res(r68_92),.clk(clk),.wout(w68_92));
	PE pe68_93(.x(x93),.w(w68_92),.acc(r68_92),.res(r68_93),.clk(clk),.wout(w68_93));
	PE pe68_94(.x(x94),.w(w68_93),.acc(r68_93),.res(r68_94),.clk(clk),.wout(w68_94));
	PE pe68_95(.x(x95),.w(w68_94),.acc(r68_94),.res(r68_95),.clk(clk),.wout(w68_95));
	PE pe68_96(.x(x96),.w(w68_95),.acc(r68_95),.res(r68_96),.clk(clk),.wout(w68_96));
	PE pe68_97(.x(x97),.w(w68_96),.acc(r68_96),.res(r68_97),.clk(clk),.wout(w68_97));
	PE pe68_98(.x(x98),.w(w68_97),.acc(r68_97),.res(r68_98),.clk(clk),.wout(w68_98));
	PE pe68_99(.x(x99),.w(w68_98),.acc(r68_98),.res(r68_99),.clk(clk),.wout(w68_99));
	PE pe68_100(.x(x100),.w(w68_99),.acc(r68_99),.res(r68_100),.clk(clk),.wout(w68_100));
	PE pe68_101(.x(x101),.w(w68_100),.acc(r68_100),.res(r68_101),.clk(clk),.wout(w68_101));
	PE pe68_102(.x(x102),.w(w68_101),.acc(r68_101),.res(r68_102),.clk(clk),.wout(w68_102));
	PE pe68_103(.x(x103),.w(w68_102),.acc(r68_102),.res(r68_103),.clk(clk),.wout(w68_103));
	PE pe68_104(.x(x104),.w(w68_103),.acc(r68_103),.res(r68_104),.clk(clk),.wout(w68_104));
	PE pe68_105(.x(x105),.w(w68_104),.acc(r68_104),.res(r68_105),.clk(clk),.wout(w68_105));
	PE pe68_106(.x(x106),.w(w68_105),.acc(r68_105),.res(r68_106),.clk(clk),.wout(w68_106));
	PE pe68_107(.x(x107),.w(w68_106),.acc(r68_106),.res(r68_107),.clk(clk),.wout(w68_107));
	PE pe68_108(.x(x108),.w(w68_107),.acc(r68_107),.res(r68_108),.clk(clk),.wout(w68_108));
	PE pe68_109(.x(x109),.w(w68_108),.acc(r68_108),.res(r68_109),.clk(clk),.wout(w68_109));
	PE pe68_110(.x(x110),.w(w68_109),.acc(r68_109),.res(r68_110),.clk(clk),.wout(w68_110));
	PE pe68_111(.x(x111),.w(w68_110),.acc(r68_110),.res(r68_111),.clk(clk),.wout(w68_111));
	PE pe68_112(.x(x112),.w(w68_111),.acc(r68_111),.res(r68_112),.clk(clk),.wout(w68_112));
	PE pe68_113(.x(x113),.w(w68_112),.acc(r68_112),.res(r68_113),.clk(clk),.wout(w68_113));
	PE pe68_114(.x(x114),.w(w68_113),.acc(r68_113),.res(r68_114),.clk(clk),.wout(w68_114));
	PE pe68_115(.x(x115),.w(w68_114),.acc(r68_114),.res(r68_115),.clk(clk),.wout(w68_115));
	PE pe68_116(.x(x116),.w(w68_115),.acc(r68_115),.res(r68_116),.clk(clk),.wout(w68_116));
	PE pe68_117(.x(x117),.w(w68_116),.acc(r68_116),.res(r68_117),.clk(clk),.wout(w68_117));
	PE pe68_118(.x(x118),.w(w68_117),.acc(r68_117),.res(r68_118),.clk(clk),.wout(w68_118));
	PE pe68_119(.x(x119),.w(w68_118),.acc(r68_118),.res(r68_119),.clk(clk),.wout(w68_119));
	PE pe68_120(.x(x120),.w(w68_119),.acc(r68_119),.res(r68_120),.clk(clk),.wout(w68_120));
	PE pe68_121(.x(x121),.w(w68_120),.acc(r68_120),.res(r68_121),.clk(clk),.wout(w68_121));
	PE pe68_122(.x(x122),.w(w68_121),.acc(r68_121),.res(r68_122),.clk(clk),.wout(w68_122));
	PE pe68_123(.x(x123),.w(w68_122),.acc(r68_122),.res(r68_123),.clk(clk),.wout(w68_123));
	PE pe68_124(.x(x124),.w(w68_123),.acc(r68_123),.res(r68_124),.clk(clk),.wout(w68_124));
	PE pe68_125(.x(x125),.w(w68_124),.acc(r68_124),.res(r68_125),.clk(clk),.wout(w68_125));
	PE pe68_126(.x(x126),.w(w68_125),.acc(r68_125),.res(r68_126),.clk(clk),.wout(w68_126));
	PE pe68_127(.x(x127),.w(w68_126),.acc(r68_126),.res(result68),.clk(clk),.wout(weight68));

	PE pe69_0(.x(x0),.w(w69),.acc(32'h0),.res(r69_0),.clk(clk),.wout(w69_0));
	PE pe69_1(.x(x1),.w(w69_0),.acc(r69_0),.res(r69_1),.clk(clk),.wout(w69_1));
	PE pe69_2(.x(x2),.w(w69_1),.acc(r69_1),.res(r69_2),.clk(clk),.wout(w69_2));
	PE pe69_3(.x(x3),.w(w69_2),.acc(r69_2),.res(r69_3),.clk(clk),.wout(w69_3));
	PE pe69_4(.x(x4),.w(w69_3),.acc(r69_3),.res(r69_4),.clk(clk),.wout(w69_4));
	PE pe69_5(.x(x5),.w(w69_4),.acc(r69_4),.res(r69_5),.clk(clk),.wout(w69_5));
	PE pe69_6(.x(x6),.w(w69_5),.acc(r69_5),.res(r69_6),.clk(clk),.wout(w69_6));
	PE pe69_7(.x(x7),.w(w69_6),.acc(r69_6),.res(r69_7),.clk(clk),.wout(w69_7));
	PE pe69_8(.x(x8),.w(w69_7),.acc(r69_7),.res(r69_8),.clk(clk),.wout(w69_8));
	PE pe69_9(.x(x9),.w(w69_8),.acc(r69_8),.res(r69_9),.clk(clk),.wout(w69_9));
	PE pe69_10(.x(x10),.w(w69_9),.acc(r69_9),.res(r69_10),.clk(clk),.wout(w69_10));
	PE pe69_11(.x(x11),.w(w69_10),.acc(r69_10),.res(r69_11),.clk(clk),.wout(w69_11));
	PE pe69_12(.x(x12),.w(w69_11),.acc(r69_11),.res(r69_12),.clk(clk),.wout(w69_12));
	PE pe69_13(.x(x13),.w(w69_12),.acc(r69_12),.res(r69_13),.clk(clk),.wout(w69_13));
	PE pe69_14(.x(x14),.w(w69_13),.acc(r69_13),.res(r69_14),.clk(clk),.wout(w69_14));
	PE pe69_15(.x(x15),.w(w69_14),.acc(r69_14),.res(r69_15),.clk(clk),.wout(w69_15));
	PE pe69_16(.x(x16),.w(w69_15),.acc(r69_15),.res(r69_16),.clk(clk),.wout(w69_16));
	PE pe69_17(.x(x17),.w(w69_16),.acc(r69_16),.res(r69_17),.clk(clk),.wout(w69_17));
	PE pe69_18(.x(x18),.w(w69_17),.acc(r69_17),.res(r69_18),.clk(clk),.wout(w69_18));
	PE pe69_19(.x(x19),.w(w69_18),.acc(r69_18),.res(r69_19),.clk(clk),.wout(w69_19));
	PE pe69_20(.x(x20),.w(w69_19),.acc(r69_19),.res(r69_20),.clk(clk),.wout(w69_20));
	PE pe69_21(.x(x21),.w(w69_20),.acc(r69_20),.res(r69_21),.clk(clk),.wout(w69_21));
	PE pe69_22(.x(x22),.w(w69_21),.acc(r69_21),.res(r69_22),.clk(clk),.wout(w69_22));
	PE pe69_23(.x(x23),.w(w69_22),.acc(r69_22),.res(r69_23),.clk(clk),.wout(w69_23));
	PE pe69_24(.x(x24),.w(w69_23),.acc(r69_23),.res(r69_24),.clk(clk),.wout(w69_24));
	PE pe69_25(.x(x25),.w(w69_24),.acc(r69_24),.res(r69_25),.clk(clk),.wout(w69_25));
	PE pe69_26(.x(x26),.w(w69_25),.acc(r69_25),.res(r69_26),.clk(clk),.wout(w69_26));
	PE pe69_27(.x(x27),.w(w69_26),.acc(r69_26),.res(r69_27),.clk(clk),.wout(w69_27));
	PE pe69_28(.x(x28),.w(w69_27),.acc(r69_27),.res(r69_28),.clk(clk),.wout(w69_28));
	PE pe69_29(.x(x29),.w(w69_28),.acc(r69_28),.res(r69_29),.clk(clk),.wout(w69_29));
	PE pe69_30(.x(x30),.w(w69_29),.acc(r69_29),.res(r69_30),.clk(clk),.wout(w69_30));
	PE pe69_31(.x(x31),.w(w69_30),.acc(r69_30),.res(r69_31),.clk(clk),.wout(w69_31));
	PE pe69_32(.x(x32),.w(w69_31),.acc(r69_31),.res(r69_32),.clk(clk),.wout(w69_32));
	PE pe69_33(.x(x33),.w(w69_32),.acc(r69_32),.res(r69_33),.clk(clk),.wout(w69_33));
	PE pe69_34(.x(x34),.w(w69_33),.acc(r69_33),.res(r69_34),.clk(clk),.wout(w69_34));
	PE pe69_35(.x(x35),.w(w69_34),.acc(r69_34),.res(r69_35),.clk(clk),.wout(w69_35));
	PE pe69_36(.x(x36),.w(w69_35),.acc(r69_35),.res(r69_36),.clk(clk),.wout(w69_36));
	PE pe69_37(.x(x37),.w(w69_36),.acc(r69_36),.res(r69_37),.clk(clk),.wout(w69_37));
	PE pe69_38(.x(x38),.w(w69_37),.acc(r69_37),.res(r69_38),.clk(clk),.wout(w69_38));
	PE pe69_39(.x(x39),.w(w69_38),.acc(r69_38),.res(r69_39),.clk(clk),.wout(w69_39));
	PE pe69_40(.x(x40),.w(w69_39),.acc(r69_39),.res(r69_40),.clk(clk),.wout(w69_40));
	PE pe69_41(.x(x41),.w(w69_40),.acc(r69_40),.res(r69_41),.clk(clk),.wout(w69_41));
	PE pe69_42(.x(x42),.w(w69_41),.acc(r69_41),.res(r69_42),.clk(clk),.wout(w69_42));
	PE pe69_43(.x(x43),.w(w69_42),.acc(r69_42),.res(r69_43),.clk(clk),.wout(w69_43));
	PE pe69_44(.x(x44),.w(w69_43),.acc(r69_43),.res(r69_44),.clk(clk),.wout(w69_44));
	PE pe69_45(.x(x45),.w(w69_44),.acc(r69_44),.res(r69_45),.clk(clk),.wout(w69_45));
	PE pe69_46(.x(x46),.w(w69_45),.acc(r69_45),.res(r69_46),.clk(clk),.wout(w69_46));
	PE pe69_47(.x(x47),.w(w69_46),.acc(r69_46),.res(r69_47),.clk(clk),.wout(w69_47));
	PE pe69_48(.x(x48),.w(w69_47),.acc(r69_47),.res(r69_48),.clk(clk),.wout(w69_48));
	PE pe69_49(.x(x49),.w(w69_48),.acc(r69_48),.res(r69_49),.clk(clk),.wout(w69_49));
	PE pe69_50(.x(x50),.w(w69_49),.acc(r69_49),.res(r69_50),.clk(clk),.wout(w69_50));
	PE pe69_51(.x(x51),.w(w69_50),.acc(r69_50),.res(r69_51),.clk(clk),.wout(w69_51));
	PE pe69_52(.x(x52),.w(w69_51),.acc(r69_51),.res(r69_52),.clk(clk),.wout(w69_52));
	PE pe69_53(.x(x53),.w(w69_52),.acc(r69_52),.res(r69_53),.clk(clk),.wout(w69_53));
	PE pe69_54(.x(x54),.w(w69_53),.acc(r69_53),.res(r69_54),.clk(clk),.wout(w69_54));
	PE pe69_55(.x(x55),.w(w69_54),.acc(r69_54),.res(r69_55),.clk(clk),.wout(w69_55));
	PE pe69_56(.x(x56),.w(w69_55),.acc(r69_55),.res(r69_56),.clk(clk),.wout(w69_56));
	PE pe69_57(.x(x57),.w(w69_56),.acc(r69_56),.res(r69_57),.clk(clk),.wout(w69_57));
	PE pe69_58(.x(x58),.w(w69_57),.acc(r69_57),.res(r69_58),.clk(clk),.wout(w69_58));
	PE pe69_59(.x(x59),.w(w69_58),.acc(r69_58),.res(r69_59),.clk(clk),.wout(w69_59));
	PE pe69_60(.x(x60),.w(w69_59),.acc(r69_59),.res(r69_60),.clk(clk),.wout(w69_60));
	PE pe69_61(.x(x61),.w(w69_60),.acc(r69_60),.res(r69_61),.clk(clk),.wout(w69_61));
	PE pe69_62(.x(x62),.w(w69_61),.acc(r69_61),.res(r69_62),.clk(clk),.wout(w69_62));
	PE pe69_63(.x(x63),.w(w69_62),.acc(r69_62),.res(r69_63),.clk(clk),.wout(w69_63));
	PE pe69_64(.x(x64),.w(w69_63),.acc(r69_63),.res(r69_64),.clk(clk),.wout(w69_64));
	PE pe69_65(.x(x65),.w(w69_64),.acc(r69_64),.res(r69_65),.clk(clk),.wout(w69_65));
	PE pe69_66(.x(x66),.w(w69_65),.acc(r69_65),.res(r69_66),.clk(clk),.wout(w69_66));
	PE pe69_67(.x(x67),.w(w69_66),.acc(r69_66),.res(r69_67),.clk(clk),.wout(w69_67));
	PE pe69_68(.x(x68),.w(w69_67),.acc(r69_67),.res(r69_68),.clk(clk),.wout(w69_68));
	PE pe69_69(.x(x69),.w(w69_68),.acc(r69_68),.res(r69_69),.clk(clk),.wout(w69_69));
	PE pe69_70(.x(x70),.w(w69_69),.acc(r69_69),.res(r69_70),.clk(clk),.wout(w69_70));
	PE pe69_71(.x(x71),.w(w69_70),.acc(r69_70),.res(r69_71),.clk(clk),.wout(w69_71));
	PE pe69_72(.x(x72),.w(w69_71),.acc(r69_71),.res(r69_72),.clk(clk),.wout(w69_72));
	PE pe69_73(.x(x73),.w(w69_72),.acc(r69_72),.res(r69_73),.clk(clk),.wout(w69_73));
	PE pe69_74(.x(x74),.w(w69_73),.acc(r69_73),.res(r69_74),.clk(clk),.wout(w69_74));
	PE pe69_75(.x(x75),.w(w69_74),.acc(r69_74),.res(r69_75),.clk(clk),.wout(w69_75));
	PE pe69_76(.x(x76),.w(w69_75),.acc(r69_75),.res(r69_76),.clk(clk),.wout(w69_76));
	PE pe69_77(.x(x77),.w(w69_76),.acc(r69_76),.res(r69_77),.clk(clk),.wout(w69_77));
	PE pe69_78(.x(x78),.w(w69_77),.acc(r69_77),.res(r69_78),.clk(clk),.wout(w69_78));
	PE pe69_79(.x(x79),.w(w69_78),.acc(r69_78),.res(r69_79),.clk(clk),.wout(w69_79));
	PE pe69_80(.x(x80),.w(w69_79),.acc(r69_79),.res(r69_80),.clk(clk),.wout(w69_80));
	PE pe69_81(.x(x81),.w(w69_80),.acc(r69_80),.res(r69_81),.clk(clk),.wout(w69_81));
	PE pe69_82(.x(x82),.w(w69_81),.acc(r69_81),.res(r69_82),.clk(clk),.wout(w69_82));
	PE pe69_83(.x(x83),.w(w69_82),.acc(r69_82),.res(r69_83),.clk(clk),.wout(w69_83));
	PE pe69_84(.x(x84),.w(w69_83),.acc(r69_83),.res(r69_84),.clk(clk),.wout(w69_84));
	PE pe69_85(.x(x85),.w(w69_84),.acc(r69_84),.res(r69_85),.clk(clk),.wout(w69_85));
	PE pe69_86(.x(x86),.w(w69_85),.acc(r69_85),.res(r69_86),.clk(clk),.wout(w69_86));
	PE pe69_87(.x(x87),.w(w69_86),.acc(r69_86),.res(r69_87),.clk(clk),.wout(w69_87));
	PE pe69_88(.x(x88),.w(w69_87),.acc(r69_87),.res(r69_88),.clk(clk),.wout(w69_88));
	PE pe69_89(.x(x89),.w(w69_88),.acc(r69_88),.res(r69_89),.clk(clk),.wout(w69_89));
	PE pe69_90(.x(x90),.w(w69_89),.acc(r69_89),.res(r69_90),.clk(clk),.wout(w69_90));
	PE pe69_91(.x(x91),.w(w69_90),.acc(r69_90),.res(r69_91),.clk(clk),.wout(w69_91));
	PE pe69_92(.x(x92),.w(w69_91),.acc(r69_91),.res(r69_92),.clk(clk),.wout(w69_92));
	PE pe69_93(.x(x93),.w(w69_92),.acc(r69_92),.res(r69_93),.clk(clk),.wout(w69_93));
	PE pe69_94(.x(x94),.w(w69_93),.acc(r69_93),.res(r69_94),.clk(clk),.wout(w69_94));
	PE pe69_95(.x(x95),.w(w69_94),.acc(r69_94),.res(r69_95),.clk(clk),.wout(w69_95));
	PE pe69_96(.x(x96),.w(w69_95),.acc(r69_95),.res(r69_96),.clk(clk),.wout(w69_96));
	PE pe69_97(.x(x97),.w(w69_96),.acc(r69_96),.res(r69_97),.clk(clk),.wout(w69_97));
	PE pe69_98(.x(x98),.w(w69_97),.acc(r69_97),.res(r69_98),.clk(clk),.wout(w69_98));
	PE pe69_99(.x(x99),.w(w69_98),.acc(r69_98),.res(r69_99),.clk(clk),.wout(w69_99));
	PE pe69_100(.x(x100),.w(w69_99),.acc(r69_99),.res(r69_100),.clk(clk),.wout(w69_100));
	PE pe69_101(.x(x101),.w(w69_100),.acc(r69_100),.res(r69_101),.clk(clk),.wout(w69_101));
	PE pe69_102(.x(x102),.w(w69_101),.acc(r69_101),.res(r69_102),.clk(clk),.wout(w69_102));
	PE pe69_103(.x(x103),.w(w69_102),.acc(r69_102),.res(r69_103),.clk(clk),.wout(w69_103));
	PE pe69_104(.x(x104),.w(w69_103),.acc(r69_103),.res(r69_104),.clk(clk),.wout(w69_104));
	PE pe69_105(.x(x105),.w(w69_104),.acc(r69_104),.res(r69_105),.clk(clk),.wout(w69_105));
	PE pe69_106(.x(x106),.w(w69_105),.acc(r69_105),.res(r69_106),.clk(clk),.wout(w69_106));
	PE pe69_107(.x(x107),.w(w69_106),.acc(r69_106),.res(r69_107),.clk(clk),.wout(w69_107));
	PE pe69_108(.x(x108),.w(w69_107),.acc(r69_107),.res(r69_108),.clk(clk),.wout(w69_108));
	PE pe69_109(.x(x109),.w(w69_108),.acc(r69_108),.res(r69_109),.clk(clk),.wout(w69_109));
	PE pe69_110(.x(x110),.w(w69_109),.acc(r69_109),.res(r69_110),.clk(clk),.wout(w69_110));
	PE pe69_111(.x(x111),.w(w69_110),.acc(r69_110),.res(r69_111),.clk(clk),.wout(w69_111));
	PE pe69_112(.x(x112),.w(w69_111),.acc(r69_111),.res(r69_112),.clk(clk),.wout(w69_112));
	PE pe69_113(.x(x113),.w(w69_112),.acc(r69_112),.res(r69_113),.clk(clk),.wout(w69_113));
	PE pe69_114(.x(x114),.w(w69_113),.acc(r69_113),.res(r69_114),.clk(clk),.wout(w69_114));
	PE pe69_115(.x(x115),.w(w69_114),.acc(r69_114),.res(r69_115),.clk(clk),.wout(w69_115));
	PE pe69_116(.x(x116),.w(w69_115),.acc(r69_115),.res(r69_116),.clk(clk),.wout(w69_116));
	PE pe69_117(.x(x117),.w(w69_116),.acc(r69_116),.res(r69_117),.clk(clk),.wout(w69_117));
	PE pe69_118(.x(x118),.w(w69_117),.acc(r69_117),.res(r69_118),.clk(clk),.wout(w69_118));
	PE pe69_119(.x(x119),.w(w69_118),.acc(r69_118),.res(r69_119),.clk(clk),.wout(w69_119));
	PE pe69_120(.x(x120),.w(w69_119),.acc(r69_119),.res(r69_120),.clk(clk),.wout(w69_120));
	PE pe69_121(.x(x121),.w(w69_120),.acc(r69_120),.res(r69_121),.clk(clk),.wout(w69_121));
	PE pe69_122(.x(x122),.w(w69_121),.acc(r69_121),.res(r69_122),.clk(clk),.wout(w69_122));
	PE pe69_123(.x(x123),.w(w69_122),.acc(r69_122),.res(r69_123),.clk(clk),.wout(w69_123));
	PE pe69_124(.x(x124),.w(w69_123),.acc(r69_123),.res(r69_124),.clk(clk),.wout(w69_124));
	PE pe69_125(.x(x125),.w(w69_124),.acc(r69_124),.res(r69_125),.clk(clk),.wout(w69_125));
	PE pe69_126(.x(x126),.w(w69_125),.acc(r69_125),.res(r69_126),.clk(clk),.wout(w69_126));
	PE pe69_127(.x(x127),.w(w69_126),.acc(r69_126),.res(result69),.clk(clk),.wout(weight69));

	PE pe70_0(.x(x0),.w(w70),.acc(32'h0),.res(r70_0),.clk(clk),.wout(w70_0));
	PE pe70_1(.x(x1),.w(w70_0),.acc(r70_0),.res(r70_1),.clk(clk),.wout(w70_1));
	PE pe70_2(.x(x2),.w(w70_1),.acc(r70_1),.res(r70_2),.clk(clk),.wout(w70_2));
	PE pe70_3(.x(x3),.w(w70_2),.acc(r70_2),.res(r70_3),.clk(clk),.wout(w70_3));
	PE pe70_4(.x(x4),.w(w70_3),.acc(r70_3),.res(r70_4),.clk(clk),.wout(w70_4));
	PE pe70_5(.x(x5),.w(w70_4),.acc(r70_4),.res(r70_5),.clk(clk),.wout(w70_5));
	PE pe70_6(.x(x6),.w(w70_5),.acc(r70_5),.res(r70_6),.clk(clk),.wout(w70_6));
	PE pe70_7(.x(x7),.w(w70_6),.acc(r70_6),.res(r70_7),.clk(clk),.wout(w70_7));
	PE pe70_8(.x(x8),.w(w70_7),.acc(r70_7),.res(r70_8),.clk(clk),.wout(w70_8));
	PE pe70_9(.x(x9),.w(w70_8),.acc(r70_8),.res(r70_9),.clk(clk),.wout(w70_9));
	PE pe70_10(.x(x10),.w(w70_9),.acc(r70_9),.res(r70_10),.clk(clk),.wout(w70_10));
	PE pe70_11(.x(x11),.w(w70_10),.acc(r70_10),.res(r70_11),.clk(clk),.wout(w70_11));
	PE pe70_12(.x(x12),.w(w70_11),.acc(r70_11),.res(r70_12),.clk(clk),.wout(w70_12));
	PE pe70_13(.x(x13),.w(w70_12),.acc(r70_12),.res(r70_13),.clk(clk),.wout(w70_13));
	PE pe70_14(.x(x14),.w(w70_13),.acc(r70_13),.res(r70_14),.clk(clk),.wout(w70_14));
	PE pe70_15(.x(x15),.w(w70_14),.acc(r70_14),.res(r70_15),.clk(clk),.wout(w70_15));
	PE pe70_16(.x(x16),.w(w70_15),.acc(r70_15),.res(r70_16),.clk(clk),.wout(w70_16));
	PE pe70_17(.x(x17),.w(w70_16),.acc(r70_16),.res(r70_17),.clk(clk),.wout(w70_17));
	PE pe70_18(.x(x18),.w(w70_17),.acc(r70_17),.res(r70_18),.clk(clk),.wout(w70_18));
	PE pe70_19(.x(x19),.w(w70_18),.acc(r70_18),.res(r70_19),.clk(clk),.wout(w70_19));
	PE pe70_20(.x(x20),.w(w70_19),.acc(r70_19),.res(r70_20),.clk(clk),.wout(w70_20));
	PE pe70_21(.x(x21),.w(w70_20),.acc(r70_20),.res(r70_21),.clk(clk),.wout(w70_21));
	PE pe70_22(.x(x22),.w(w70_21),.acc(r70_21),.res(r70_22),.clk(clk),.wout(w70_22));
	PE pe70_23(.x(x23),.w(w70_22),.acc(r70_22),.res(r70_23),.clk(clk),.wout(w70_23));
	PE pe70_24(.x(x24),.w(w70_23),.acc(r70_23),.res(r70_24),.clk(clk),.wout(w70_24));
	PE pe70_25(.x(x25),.w(w70_24),.acc(r70_24),.res(r70_25),.clk(clk),.wout(w70_25));
	PE pe70_26(.x(x26),.w(w70_25),.acc(r70_25),.res(r70_26),.clk(clk),.wout(w70_26));
	PE pe70_27(.x(x27),.w(w70_26),.acc(r70_26),.res(r70_27),.clk(clk),.wout(w70_27));
	PE pe70_28(.x(x28),.w(w70_27),.acc(r70_27),.res(r70_28),.clk(clk),.wout(w70_28));
	PE pe70_29(.x(x29),.w(w70_28),.acc(r70_28),.res(r70_29),.clk(clk),.wout(w70_29));
	PE pe70_30(.x(x30),.w(w70_29),.acc(r70_29),.res(r70_30),.clk(clk),.wout(w70_30));
	PE pe70_31(.x(x31),.w(w70_30),.acc(r70_30),.res(r70_31),.clk(clk),.wout(w70_31));
	PE pe70_32(.x(x32),.w(w70_31),.acc(r70_31),.res(r70_32),.clk(clk),.wout(w70_32));
	PE pe70_33(.x(x33),.w(w70_32),.acc(r70_32),.res(r70_33),.clk(clk),.wout(w70_33));
	PE pe70_34(.x(x34),.w(w70_33),.acc(r70_33),.res(r70_34),.clk(clk),.wout(w70_34));
	PE pe70_35(.x(x35),.w(w70_34),.acc(r70_34),.res(r70_35),.clk(clk),.wout(w70_35));
	PE pe70_36(.x(x36),.w(w70_35),.acc(r70_35),.res(r70_36),.clk(clk),.wout(w70_36));
	PE pe70_37(.x(x37),.w(w70_36),.acc(r70_36),.res(r70_37),.clk(clk),.wout(w70_37));
	PE pe70_38(.x(x38),.w(w70_37),.acc(r70_37),.res(r70_38),.clk(clk),.wout(w70_38));
	PE pe70_39(.x(x39),.w(w70_38),.acc(r70_38),.res(r70_39),.clk(clk),.wout(w70_39));
	PE pe70_40(.x(x40),.w(w70_39),.acc(r70_39),.res(r70_40),.clk(clk),.wout(w70_40));
	PE pe70_41(.x(x41),.w(w70_40),.acc(r70_40),.res(r70_41),.clk(clk),.wout(w70_41));
	PE pe70_42(.x(x42),.w(w70_41),.acc(r70_41),.res(r70_42),.clk(clk),.wout(w70_42));
	PE pe70_43(.x(x43),.w(w70_42),.acc(r70_42),.res(r70_43),.clk(clk),.wout(w70_43));
	PE pe70_44(.x(x44),.w(w70_43),.acc(r70_43),.res(r70_44),.clk(clk),.wout(w70_44));
	PE pe70_45(.x(x45),.w(w70_44),.acc(r70_44),.res(r70_45),.clk(clk),.wout(w70_45));
	PE pe70_46(.x(x46),.w(w70_45),.acc(r70_45),.res(r70_46),.clk(clk),.wout(w70_46));
	PE pe70_47(.x(x47),.w(w70_46),.acc(r70_46),.res(r70_47),.clk(clk),.wout(w70_47));
	PE pe70_48(.x(x48),.w(w70_47),.acc(r70_47),.res(r70_48),.clk(clk),.wout(w70_48));
	PE pe70_49(.x(x49),.w(w70_48),.acc(r70_48),.res(r70_49),.clk(clk),.wout(w70_49));
	PE pe70_50(.x(x50),.w(w70_49),.acc(r70_49),.res(r70_50),.clk(clk),.wout(w70_50));
	PE pe70_51(.x(x51),.w(w70_50),.acc(r70_50),.res(r70_51),.clk(clk),.wout(w70_51));
	PE pe70_52(.x(x52),.w(w70_51),.acc(r70_51),.res(r70_52),.clk(clk),.wout(w70_52));
	PE pe70_53(.x(x53),.w(w70_52),.acc(r70_52),.res(r70_53),.clk(clk),.wout(w70_53));
	PE pe70_54(.x(x54),.w(w70_53),.acc(r70_53),.res(r70_54),.clk(clk),.wout(w70_54));
	PE pe70_55(.x(x55),.w(w70_54),.acc(r70_54),.res(r70_55),.clk(clk),.wout(w70_55));
	PE pe70_56(.x(x56),.w(w70_55),.acc(r70_55),.res(r70_56),.clk(clk),.wout(w70_56));
	PE pe70_57(.x(x57),.w(w70_56),.acc(r70_56),.res(r70_57),.clk(clk),.wout(w70_57));
	PE pe70_58(.x(x58),.w(w70_57),.acc(r70_57),.res(r70_58),.clk(clk),.wout(w70_58));
	PE pe70_59(.x(x59),.w(w70_58),.acc(r70_58),.res(r70_59),.clk(clk),.wout(w70_59));
	PE pe70_60(.x(x60),.w(w70_59),.acc(r70_59),.res(r70_60),.clk(clk),.wout(w70_60));
	PE pe70_61(.x(x61),.w(w70_60),.acc(r70_60),.res(r70_61),.clk(clk),.wout(w70_61));
	PE pe70_62(.x(x62),.w(w70_61),.acc(r70_61),.res(r70_62),.clk(clk),.wout(w70_62));
	PE pe70_63(.x(x63),.w(w70_62),.acc(r70_62),.res(r70_63),.clk(clk),.wout(w70_63));
	PE pe70_64(.x(x64),.w(w70_63),.acc(r70_63),.res(r70_64),.clk(clk),.wout(w70_64));
	PE pe70_65(.x(x65),.w(w70_64),.acc(r70_64),.res(r70_65),.clk(clk),.wout(w70_65));
	PE pe70_66(.x(x66),.w(w70_65),.acc(r70_65),.res(r70_66),.clk(clk),.wout(w70_66));
	PE pe70_67(.x(x67),.w(w70_66),.acc(r70_66),.res(r70_67),.clk(clk),.wout(w70_67));
	PE pe70_68(.x(x68),.w(w70_67),.acc(r70_67),.res(r70_68),.clk(clk),.wout(w70_68));
	PE pe70_69(.x(x69),.w(w70_68),.acc(r70_68),.res(r70_69),.clk(clk),.wout(w70_69));
	PE pe70_70(.x(x70),.w(w70_69),.acc(r70_69),.res(r70_70),.clk(clk),.wout(w70_70));
	PE pe70_71(.x(x71),.w(w70_70),.acc(r70_70),.res(r70_71),.clk(clk),.wout(w70_71));
	PE pe70_72(.x(x72),.w(w70_71),.acc(r70_71),.res(r70_72),.clk(clk),.wout(w70_72));
	PE pe70_73(.x(x73),.w(w70_72),.acc(r70_72),.res(r70_73),.clk(clk),.wout(w70_73));
	PE pe70_74(.x(x74),.w(w70_73),.acc(r70_73),.res(r70_74),.clk(clk),.wout(w70_74));
	PE pe70_75(.x(x75),.w(w70_74),.acc(r70_74),.res(r70_75),.clk(clk),.wout(w70_75));
	PE pe70_76(.x(x76),.w(w70_75),.acc(r70_75),.res(r70_76),.clk(clk),.wout(w70_76));
	PE pe70_77(.x(x77),.w(w70_76),.acc(r70_76),.res(r70_77),.clk(clk),.wout(w70_77));
	PE pe70_78(.x(x78),.w(w70_77),.acc(r70_77),.res(r70_78),.clk(clk),.wout(w70_78));
	PE pe70_79(.x(x79),.w(w70_78),.acc(r70_78),.res(r70_79),.clk(clk),.wout(w70_79));
	PE pe70_80(.x(x80),.w(w70_79),.acc(r70_79),.res(r70_80),.clk(clk),.wout(w70_80));
	PE pe70_81(.x(x81),.w(w70_80),.acc(r70_80),.res(r70_81),.clk(clk),.wout(w70_81));
	PE pe70_82(.x(x82),.w(w70_81),.acc(r70_81),.res(r70_82),.clk(clk),.wout(w70_82));
	PE pe70_83(.x(x83),.w(w70_82),.acc(r70_82),.res(r70_83),.clk(clk),.wout(w70_83));
	PE pe70_84(.x(x84),.w(w70_83),.acc(r70_83),.res(r70_84),.clk(clk),.wout(w70_84));
	PE pe70_85(.x(x85),.w(w70_84),.acc(r70_84),.res(r70_85),.clk(clk),.wout(w70_85));
	PE pe70_86(.x(x86),.w(w70_85),.acc(r70_85),.res(r70_86),.clk(clk),.wout(w70_86));
	PE pe70_87(.x(x87),.w(w70_86),.acc(r70_86),.res(r70_87),.clk(clk),.wout(w70_87));
	PE pe70_88(.x(x88),.w(w70_87),.acc(r70_87),.res(r70_88),.clk(clk),.wout(w70_88));
	PE pe70_89(.x(x89),.w(w70_88),.acc(r70_88),.res(r70_89),.clk(clk),.wout(w70_89));
	PE pe70_90(.x(x90),.w(w70_89),.acc(r70_89),.res(r70_90),.clk(clk),.wout(w70_90));
	PE pe70_91(.x(x91),.w(w70_90),.acc(r70_90),.res(r70_91),.clk(clk),.wout(w70_91));
	PE pe70_92(.x(x92),.w(w70_91),.acc(r70_91),.res(r70_92),.clk(clk),.wout(w70_92));
	PE pe70_93(.x(x93),.w(w70_92),.acc(r70_92),.res(r70_93),.clk(clk),.wout(w70_93));
	PE pe70_94(.x(x94),.w(w70_93),.acc(r70_93),.res(r70_94),.clk(clk),.wout(w70_94));
	PE pe70_95(.x(x95),.w(w70_94),.acc(r70_94),.res(r70_95),.clk(clk),.wout(w70_95));
	PE pe70_96(.x(x96),.w(w70_95),.acc(r70_95),.res(r70_96),.clk(clk),.wout(w70_96));
	PE pe70_97(.x(x97),.w(w70_96),.acc(r70_96),.res(r70_97),.clk(clk),.wout(w70_97));
	PE pe70_98(.x(x98),.w(w70_97),.acc(r70_97),.res(r70_98),.clk(clk),.wout(w70_98));
	PE pe70_99(.x(x99),.w(w70_98),.acc(r70_98),.res(r70_99),.clk(clk),.wout(w70_99));
	PE pe70_100(.x(x100),.w(w70_99),.acc(r70_99),.res(r70_100),.clk(clk),.wout(w70_100));
	PE pe70_101(.x(x101),.w(w70_100),.acc(r70_100),.res(r70_101),.clk(clk),.wout(w70_101));
	PE pe70_102(.x(x102),.w(w70_101),.acc(r70_101),.res(r70_102),.clk(clk),.wout(w70_102));
	PE pe70_103(.x(x103),.w(w70_102),.acc(r70_102),.res(r70_103),.clk(clk),.wout(w70_103));
	PE pe70_104(.x(x104),.w(w70_103),.acc(r70_103),.res(r70_104),.clk(clk),.wout(w70_104));
	PE pe70_105(.x(x105),.w(w70_104),.acc(r70_104),.res(r70_105),.clk(clk),.wout(w70_105));
	PE pe70_106(.x(x106),.w(w70_105),.acc(r70_105),.res(r70_106),.clk(clk),.wout(w70_106));
	PE pe70_107(.x(x107),.w(w70_106),.acc(r70_106),.res(r70_107),.clk(clk),.wout(w70_107));
	PE pe70_108(.x(x108),.w(w70_107),.acc(r70_107),.res(r70_108),.clk(clk),.wout(w70_108));
	PE pe70_109(.x(x109),.w(w70_108),.acc(r70_108),.res(r70_109),.clk(clk),.wout(w70_109));
	PE pe70_110(.x(x110),.w(w70_109),.acc(r70_109),.res(r70_110),.clk(clk),.wout(w70_110));
	PE pe70_111(.x(x111),.w(w70_110),.acc(r70_110),.res(r70_111),.clk(clk),.wout(w70_111));
	PE pe70_112(.x(x112),.w(w70_111),.acc(r70_111),.res(r70_112),.clk(clk),.wout(w70_112));
	PE pe70_113(.x(x113),.w(w70_112),.acc(r70_112),.res(r70_113),.clk(clk),.wout(w70_113));
	PE pe70_114(.x(x114),.w(w70_113),.acc(r70_113),.res(r70_114),.clk(clk),.wout(w70_114));
	PE pe70_115(.x(x115),.w(w70_114),.acc(r70_114),.res(r70_115),.clk(clk),.wout(w70_115));
	PE pe70_116(.x(x116),.w(w70_115),.acc(r70_115),.res(r70_116),.clk(clk),.wout(w70_116));
	PE pe70_117(.x(x117),.w(w70_116),.acc(r70_116),.res(r70_117),.clk(clk),.wout(w70_117));
	PE pe70_118(.x(x118),.w(w70_117),.acc(r70_117),.res(r70_118),.clk(clk),.wout(w70_118));
	PE pe70_119(.x(x119),.w(w70_118),.acc(r70_118),.res(r70_119),.clk(clk),.wout(w70_119));
	PE pe70_120(.x(x120),.w(w70_119),.acc(r70_119),.res(r70_120),.clk(clk),.wout(w70_120));
	PE pe70_121(.x(x121),.w(w70_120),.acc(r70_120),.res(r70_121),.clk(clk),.wout(w70_121));
	PE pe70_122(.x(x122),.w(w70_121),.acc(r70_121),.res(r70_122),.clk(clk),.wout(w70_122));
	PE pe70_123(.x(x123),.w(w70_122),.acc(r70_122),.res(r70_123),.clk(clk),.wout(w70_123));
	PE pe70_124(.x(x124),.w(w70_123),.acc(r70_123),.res(r70_124),.clk(clk),.wout(w70_124));
	PE pe70_125(.x(x125),.w(w70_124),.acc(r70_124),.res(r70_125),.clk(clk),.wout(w70_125));
	PE pe70_126(.x(x126),.w(w70_125),.acc(r70_125),.res(r70_126),.clk(clk),.wout(w70_126));
	PE pe70_127(.x(x127),.w(w70_126),.acc(r70_126),.res(result70),.clk(clk),.wout(weight70));

	PE pe71_0(.x(x0),.w(w71),.acc(32'h0),.res(r71_0),.clk(clk),.wout(w71_0));
	PE pe71_1(.x(x1),.w(w71_0),.acc(r71_0),.res(r71_1),.clk(clk),.wout(w71_1));
	PE pe71_2(.x(x2),.w(w71_1),.acc(r71_1),.res(r71_2),.clk(clk),.wout(w71_2));
	PE pe71_3(.x(x3),.w(w71_2),.acc(r71_2),.res(r71_3),.clk(clk),.wout(w71_3));
	PE pe71_4(.x(x4),.w(w71_3),.acc(r71_3),.res(r71_4),.clk(clk),.wout(w71_4));
	PE pe71_5(.x(x5),.w(w71_4),.acc(r71_4),.res(r71_5),.clk(clk),.wout(w71_5));
	PE pe71_6(.x(x6),.w(w71_5),.acc(r71_5),.res(r71_6),.clk(clk),.wout(w71_6));
	PE pe71_7(.x(x7),.w(w71_6),.acc(r71_6),.res(r71_7),.clk(clk),.wout(w71_7));
	PE pe71_8(.x(x8),.w(w71_7),.acc(r71_7),.res(r71_8),.clk(clk),.wout(w71_8));
	PE pe71_9(.x(x9),.w(w71_8),.acc(r71_8),.res(r71_9),.clk(clk),.wout(w71_9));
	PE pe71_10(.x(x10),.w(w71_9),.acc(r71_9),.res(r71_10),.clk(clk),.wout(w71_10));
	PE pe71_11(.x(x11),.w(w71_10),.acc(r71_10),.res(r71_11),.clk(clk),.wout(w71_11));
	PE pe71_12(.x(x12),.w(w71_11),.acc(r71_11),.res(r71_12),.clk(clk),.wout(w71_12));
	PE pe71_13(.x(x13),.w(w71_12),.acc(r71_12),.res(r71_13),.clk(clk),.wout(w71_13));
	PE pe71_14(.x(x14),.w(w71_13),.acc(r71_13),.res(r71_14),.clk(clk),.wout(w71_14));
	PE pe71_15(.x(x15),.w(w71_14),.acc(r71_14),.res(r71_15),.clk(clk),.wout(w71_15));
	PE pe71_16(.x(x16),.w(w71_15),.acc(r71_15),.res(r71_16),.clk(clk),.wout(w71_16));
	PE pe71_17(.x(x17),.w(w71_16),.acc(r71_16),.res(r71_17),.clk(clk),.wout(w71_17));
	PE pe71_18(.x(x18),.w(w71_17),.acc(r71_17),.res(r71_18),.clk(clk),.wout(w71_18));
	PE pe71_19(.x(x19),.w(w71_18),.acc(r71_18),.res(r71_19),.clk(clk),.wout(w71_19));
	PE pe71_20(.x(x20),.w(w71_19),.acc(r71_19),.res(r71_20),.clk(clk),.wout(w71_20));
	PE pe71_21(.x(x21),.w(w71_20),.acc(r71_20),.res(r71_21),.clk(clk),.wout(w71_21));
	PE pe71_22(.x(x22),.w(w71_21),.acc(r71_21),.res(r71_22),.clk(clk),.wout(w71_22));
	PE pe71_23(.x(x23),.w(w71_22),.acc(r71_22),.res(r71_23),.clk(clk),.wout(w71_23));
	PE pe71_24(.x(x24),.w(w71_23),.acc(r71_23),.res(r71_24),.clk(clk),.wout(w71_24));
	PE pe71_25(.x(x25),.w(w71_24),.acc(r71_24),.res(r71_25),.clk(clk),.wout(w71_25));
	PE pe71_26(.x(x26),.w(w71_25),.acc(r71_25),.res(r71_26),.clk(clk),.wout(w71_26));
	PE pe71_27(.x(x27),.w(w71_26),.acc(r71_26),.res(r71_27),.clk(clk),.wout(w71_27));
	PE pe71_28(.x(x28),.w(w71_27),.acc(r71_27),.res(r71_28),.clk(clk),.wout(w71_28));
	PE pe71_29(.x(x29),.w(w71_28),.acc(r71_28),.res(r71_29),.clk(clk),.wout(w71_29));
	PE pe71_30(.x(x30),.w(w71_29),.acc(r71_29),.res(r71_30),.clk(clk),.wout(w71_30));
	PE pe71_31(.x(x31),.w(w71_30),.acc(r71_30),.res(r71_31),.clk(clk),.wout(w71_31));
	PE pe71_32(.x(x32),.w(w71_31),.acc(r71_31),.res(r71_32),.clk(clk),.wout(w71_32));
	PE pe71_33(.x(x33),.w(w71_32),.acc(r71_32),.res(r71_33),.clk(clk),.wout(w71_33));
	PE pe71_34(.x(x34),.w(w71_33),.acc(r71_33),.res(r71_34),.clk(clk),.wout(w71_34));
	PE pe71_35(.x(x35),.w(w71_34),.acc(r71_34),.res(r71_35),.clk(clk),.wout(w71_35));
	PE pe71_36(.x(x36),.w(w71_35),.acc(r71_35),.res(r71_36),.clk(clk),.wout(w71_36));
	PE pe71_37(.x(x37),.w(w71_36),.acc(r71_36),.res(r71_37),.clk(clk),.wout(w71_37));
	PE pe71_38(.x(x38),.w(w71_37),.acc(r71_37),.res(r71_38),.clk(clk),.wout(w71_38));
	PE pe71_39(.x(x39),.w(w71_38),.acc(r71_38),.res(r71_39),.clk(clk),.wout(w71_39));
	PE pe71_40(.x(x40),.w(w71_39),.acc(r71_39),.res(r71_40),.clk(clk),.wout(w71_40));
	PE pe71_41(.x(x41),.w(w71_40),.acc(r71_40),.res(r71_41),.clk(clk),.wout(w71_41));
	PE pe71_42(.x(x42),.w(w71_41),.acc(r71_41),.res(r71_42),.clk(clk),.wout(w71_42));
	PE pe71_43(.x(x43),.w(w71_42),.acc(r71_42),.res(r71_43),.clk(clk),.wout(w71_43));
	PE pe71_44(.x(x44),.w(w71_43),.acc(r71_43),.res(r71_44),.clk(clk),.wout(w71_44));
	PE pe71_45(.x(x45),.w(w71_44),.acc(r71_44),.res(r71_45),.clk(clk),.wout(w71_45));
	PE pe71_46(.x(x46),.w(w71_45),.acc(r71_45),.res(r71_46),.clk(clk),.wout(w71_46));
	PE pe71_47(.x(x47),.w(w71_46),.acc(r71_46),.res(r71_47),.clk(clk),.wout(w71_47));
	PE pe71_48(.x(x48),.w(w71_47),.acc(r71_47),.res(r71_48),.clk(clk),.wout(w71_48));
	PE pe71_49(.x(x49),.w(w71_48),.acc(r71_48),.res(r71_49),.clk(clk),.wout(w71_49));
	PE pe71_50(.x(x50),.w(w71_49),.acc(r71_49),.res(r71_50),.clk(clk),.wout(w71_50));
	PE pe71_51(.x(x51),.w(w71_50),.acc(r71_50),.res(r71_51),.clk(clk),.wout(w71_51));
	PE pe71_52(.x(x52),.w(w71_51),.acc(r71_51),.res(r71_52),.clk(clk),.wout(w71_52));
	PE pe71_53(.x(x53),.w(w71_52),.acc(r71_52),.res(r71_53),.clk(clk),.wout(w71_53));
	PE pe71_54(.x(x54),.w(w71_53),.acc(r71_53),.res(r71_54),.clk(clk),.wout(w71_54));
	PE pe71_55(.x(x55),.w(w71_54),.acc(r71_54),.res(r71_55),.clk(clk),.wout(w71_55));
	PE pe71_56(.x(x56),.w(w71_55),.acc(r71_55),.res(r71_56),.clk(clk),.wout(w71_56));
	PE pe71_57(.x(x57),.w(w71_56),.acc(r71_56),.res(r71_57),.clk(clk),.wout(w71_57));
	PE pe71_58(.x(x58),.w(w71_57),.acc(r71_57),.res(r71_58),.clk(clk),.wout(w71_58));
	PE pe71_59(.x(x59),.w(w71_58),.acc(r71_58),.res(r71_59),.clk(clk),.wout(w71_59));
	PE pe71_60(.x(x60),.w(w71_59),.acc(r71_59),.res(r71_60),.clk(clk),.wout(w71_60));
	PE pe71_61(.x(x61),.w(w71_60),.acc(r71_60),.res(r71_61),.clk(clk),.wout(w71_61));
	PE pe71_62(.x(x62),.w(w71_61),.acc(r71_61),.res(r71_62),.clk(clk),.wout(w71_62));
	PE pe71_63(.x(x63),.w(w71_62),.acc(r71_62),.res(r71_63),.clk(clk),.wout(w71_63));
	PE pe71_64(.x(x64),.w(w71_63),.acc(r71_63),.res(r71_64),.clk(clk),.wout(w71_64));
	PE pe71_65(.x(x65),.w(w71_64),.acc(r71_64),.res(r71_65),.clk(clk),.wout(w71_65));
	PE pe71_66(.x(x66),.w(w71_65),.acc(r71_65),.res(r71_66),.clk(clk),.wout(w71_66));
	PE pe71_67(.x(x67),.w(w71_66),.acc(r71_66),.res(r71_67),.clk(clk),.wout(w71_67));
	PE pe71_68(.x(x68),.w(w71_67),.acc(r71_67),.res(r71_68),.clk(clk),.wout(w71_68));
	PE pe71_69(.x(x69),.w(w71_68),.acc(r71_68),.res(r71_69),.clk(clk),.wout(w71_69));
	PE pe71_70(.x(x70),.w(w71_69),.acc(r71_69),.res(r71_70),.clk(clk),.wout(w71_70));
	PE pe71_71(.x(x71),.w(w71_70),.acc(r71_70),.res(r71_71),.clk(clk),.wout(w71_71));
	PE pe71_72(.x(x72),.w(w71_71),.acc(r71_71),.res(r71_72),.clk(clk),.wout(w71_72));
	PE pe71_73(.x(x73),.w(w71_72),.acc(r71_72),.res(r71_73),.clk(clk),.wout(w71_73));
	PE pe71_74(.x(x74),.w(w71_73),.acc(r71_73),.res(r71_74),.clk(clk),.wout(w71_74));
	PE pe71_75(.x(x75),.w(w71_74),.acc(r71_74),.res(r71_75),.clk(clk),.wout(w71_75));
	PE pe71_76(.x(x76),.w(w71_75),.acc(r71_75),.res(r71_76),.clk(clk),.wout(w71_76));
	PE pe71_77(.x(x77),.w(w71_76),.acc(r71_76),.res(r71_77),.clk(clk),.wout(w71_77));
	PE pe71_78(.x(x78),.w(w71_77),.acc(r71_77),.res(r71_78),.clk(clk),.wout(w71_78));
	PE pe71_79(.x(x79),.w(w71_78),.acc(r71_78),.res(r71_79),.clk(clk),.wout(w71_79));
	PE pe71_80(.x(x80),.w(w71_79),.acc(r71_79),.res(r71_80),.clk(clk),.wout(w71_80));
	PE pe71_81(.x(x81),.w(w71_80),.acc(r71_80),.res(r71_81),.clk(clk),.wout(w71_81));
	PE pe71_82(.x(x82),.w(w71_81),.acc(r71_81),.res(r71_82),.clk(clk),.wout(w71_82));
	PE pe71_83(.x(x83),.w(w71_82),.acc(r71_82),.res(r71_83),.clk(clk),.wout(w71_83));
	PE pe71_84(.x(x84),.w(w71_83),.acc(r71_83),.res(r71_84),.clk(clk),.wout(w71_84));
	PE pe71_85(.x(x85),.w(w71_84),.acc(r71_84),.res(r71_85),.clk(clk),.wout(w71_85));
	PE pe71_86(.x(x86),.w(w71_85),.acc(r71_85),.res(r71_86),.clk(clk),.wout(w71_86));
	PE pe71_87(.x(x87),.w(w71_86),.acc(r71_86),.res(r71_87),.clk(clk),.wout(w71_87));
	PE pe71_88(.x(x88),.w(w71_87),.acc(r71_87),.res(r71_88),.clk(clk),.wout(w71_88));
	PE pe71_89(.x(x89),.w(w71_88),.acc(r71_88),.res(r71_89),.clk(clk),.wout(w71_89));
	PE pe71_90(.x(x90),.w(w71_89),.acc(r71_89),.res(r71_90),.clk(clk),.wout(w71_90));
	PE pe71_91(.x(x91),.w(w71_90),.acc(r71_90),.res(r71_91),.clk(clk),.wout(w71_91));
	PE pe71_92(.x(x92),.w(w71_91),.acc(r71_91),.res(r71_92),.clk(clk),.wout(w71_92));
	PE pe71_93(.x(x93),.w(w71_92),.acc(r71_92),.res(r71_93),.clk(clk),.wout(w71_93));
	PE pe71_94(.x(x94),.w(w71_93),.acc(r71_93),.res(r71_94),.clk(clk),.wout(w71_94));
	PE pe71_95(.x(x95),.w(w71_94),.acc(r71_94),.res(r71_95),.clk(clk),.wout(w71_95));
	PE pe71_96(.x(x96),.w(w71_95),.acc(r71_95),.res(r71_96),.clk(clk),.wout(w71_96));
	PE pe71_97(.x(x97),.w(w71_96),.acc(r71_96),.res(r71_97),.clk(clk),.wout(w71_97));
	PE pe71_98(.x(x98),.w(w71_97),.acc(r71_97),.res(r71_98),.clk(clk),.wout(w71_98));
	PE pe71_99(.x(x99),.w(w71_98),.acc(r71_98),.res(r71_99),.clk(clk),.wout(w71_99));
	PE pe71_100(.x(x100),.w(w71_99),.acc(r71_99),.res(r71_100),.clk(clk),.wout(w71_100));
	PE pe71_101(.x(x101),.w(w71_100),.acc(r71_100),.res(r71_101),.clk(clk),.wout(w71_101));
	PE pe71_102(.x(x102),.w(w71_101),.acc(r71_101),.res(r71_102),.clk(clk),.wout(w71_102));
	PE pe71_103(.x(x103),.w(w71_102),.acc(r71_102),.res(r71_103),.clk(clk),.wout(w71_103));
	PE pe71_104(.x(x104),.w(w71_103),.acc(r71_103),.res(r71_104),.clk(clk),.wout(w71_104));
	PE pe71_105(.x(x105),.w(w71_104),.acc(r71_104),.res(r71_105),.clk(clk),.wout(w71_105));
	PE pe71_106(.x(x106),.w(w71_105),.acc(r71_105),.res(r71_106),.clk(clk),.wout(w71_106));
	PE pe71_107(.x(x107),.w(w71_106),.acc(r71_106),.res(r71_107),.clk(clk),.wout(w71_107));
	PE pe71_108(.x(x108),.w(w71_107),.acc(r71_107),.res(r71_108),.clk(clk),.wout(w71_108));
	PE pe71_109(.x(x109),.w(w71_108),.acc(r71_108),.res(r71_109),.clk(clk),.wout(w71_109));
	PE pe71_110(.x(x110),.w(w71_109),.acc(r71_109),.res(r71_110),.clk(clk),.wout(w71_110));
	PE pe71_111(.x(x111),.w(w71_110),.acc(r71_110),.res(r71_111),.clk(clk),.wout(w71_111));
	PE pe71_112(.x(x112),.w(w71_111),.acc(r71_111),.res(r71_112),.clk(clk),.wout(w71_112));
	PE pe71_113(.x(x113),.w(w71_112),.acc(r71_112),.res(r71_113),.clk(clk),.wout(w71_113));
	PE pe71_114(.x(x114),.w(w71_113),.acc(r71_113),.res(r71_114),.clk(clk),.wout(w71_114));
	PE pe71_115(.x(x115),.w(w71_114),.acc(r71_114),.res(r71_115),.clk(clk),.wout(w71_115));
	PE pe71_116(.x(x116),.w(w71_115),.acc(r71_115),.res(r71_116),.clk(clk),.wout(w71_116));
	PE pe71_117(.x(x117),.w(w71_116),.acc(r71_116),.res(r71_117),.clk(clk),.wout(w71_117));
	PE pe71_118(.x(x118),.w(w71_117),.acc(r71_117),.res(r71_118),.clk(clk),.wout(w71_118));
	PE pe71_119(.x(x119),.w(w71_118),.acc(r71_118),.res(r71_119),.clk(clk),.wout(w71_119));
	PE pe71_120(.x(x120),.w(w71_119),.acc(r71_119),.res(r71_120),.clk(clk),.wout(w71_120));
	PE pe71_121(.x(x121),.w(w71_120),.acc(r71_120),.res(r71_121),.clk(clk),.wout(w71_121));
	PE pe71_122(.x(x122),.w(w71_121),.acc(r71_121),.res(r71_122),.clk(clk),.wout(w71_122));
	PE pe71_123(.x(x123),.w(w71_122),.acc(r71_122),.res(r71_123),.clk(clk),.wout(w71_123));
	PE pe71_124(.x(x124),.w(w71_123),.acc(r71_123),.res(r71_124),.clk(clk),.wout(w71_124));
	PE pe71_125(.x(x125),.w(w71_124),.acc(r71_124),.res(r71_125),.clk(clk),.wout(w71_125));
	PE pe71_126(.x(x126),.w(w71_125),.acc(r71_125),.res(r71_126),.clk(clk),.wout(w71_126));
	PE pe71_127(.x(x127),.w(w71_126),.acc(r71_126),.res(result71),.clk(clk),.wout(weight71));

	PE pe72_0(.x(x0),.w(w72),.acc(32'h0),.res(r72_0),.clk(clk),.wout(w72_0));
	PE pe72_1(.x(x1),.w(w72_0),.acc(r72_0),.res(r72_1),.clk(clk),.wout(w72_1));
	PE pe72_2(.x(x2),.w(w72_1),.acc(r72_1),.res(r72_2),.clk(clk),.wout(w72_2));
	PE pe72_3(.x(x3),.w(w72_2),.acc(r72_2),.res(r72_3),.clk(clk),.wout(w72_3));
	PE pe72_4(.x(x4),.w(w72_3),.acc(r72_3),.res(r72_4),.clk(clk),.wout(w72_4));
	PE pe72_5(.x(x5),.w(w72_4),.acc(r72_4),.res(r72_5),.clk(clk),.wout(w72_5));
	PE pe72_6(.x(x6),.w(w72_5),.acc(r72_5),.res(r72_6),.clk(clk),.wout(w72_6));
	PE pe72_7(.x(x7),.w(w72_6),.acc(r72_6),.res(r72_7),.clk(clk),.wout(w72_7));
	PE pe72_8(.x(x8),.w(w72_7),.acc(r72_7),.res(r72_8),.clk(clk),.wout(w72_8));
	PE pe72_9(.x(x9),.w(w72_8),.acc(r72_8),.res(r72_9),.clk(clk),.wout(w72_9));
	PE pe72_10(.x(x10),.w(w72_9),.acc(r72_9),.res(r72_10),.clk(clk),.wout(w72_10));
	PE pe72_11(.x(x11),.w(w72_10),.acc(r72_10),.res(r72_11),.clk(clk),.wout(w72_11));
	PE pe72_12(.x(x12),.w(w72_11),.acc(r72_11),.res(r72_12),.clk(clk),.wout(w72_12));
	PE pe72_13(.x(x13),.w(w72_12),.acc(r72_12),.res(r72_13),.clk(clk),.wout(w72_13));
	PE pe72_14(.x(x14),.w(w72_13),.acc(r72_13),.res(r72_14),.clk(clk),.wout(w72_14));
	PE pe72_15(.x(x15),.w(w72_14),.acc(r72_14),.res(r72_15),.clk(clk),.wout(w72_15));
	PE pe72_16(.x(x16),.w(w72_15),.acc(r72_15),.res(r72_16),.clk(clk),.wout(w72_16));
	PE pe72_17(.x(x17),.w(w72_16),.acc(r72_16),.res(r72_17),.clk(clk),.wout(w72_17));
	PE pe72_18(.x(x18),.w(w72_17),.acc(r72_17),.res(r72_18),.clk(clk),.wout(w72_18));
	PE pe72_19(.x(x19),.w(w72_18),.acc(r72_18),.res(r72_19),.clk(clk),.wout(w72_19));
	PE pe72_20(.x(x20),.w(w72_19),.acc(r72_19),.res(r72_20),.clk(clk),.wout(w72_20));
	PE pe72_21(.x(x21),.w(w72_20),.acc(r72_20),.res(r72_21),.clk(clk),.wout(w72_21));
	PE pe72_22(.x(x22),.w(w72_21),.acc(r72_21),.res(r72_22),.clk(clk),.wout(w72_22));
	PE pe72_23(.x(x23),.w(w72_22),.acc(r72_22),.res(r72_23),.clk(clk),.wout(w72_23));
	PE pe72_24(.x(x24),.w(w72_23),.acc(r72_23),.res(r72_24),.clk(clk),.wout(w72_24));
	PE pe72_25(.x(x25),.w(w72_24),.acc(r72_24),.res(r72_25),.clk(clk),.wout(w72_25));
	PE pe72_26(.x(x26),.w(w72_25),.acc(r72_25),.res(r72_26),.clk(clk),.wout(w72_26));
	PE pe72_27(.x(x27),.w(w72_26),.acc(r72_26),.res(r72_27),.clk(clk),.wout(w72_27));
	PE pe72_28(.x(x28),.w(w72_27),.acc(r72_27),.res(r72_28),.clk(clk),.wout(w72_28));
	PE pe72_29(.x(x29),.w(w72_28),.acc(r72_28),.res(r72_29),.clk(clk),.wout(w72_29));
	PE pe72_30(.x(x30),.w(w72_29),.acc(r72_29),.res(r72_30),.clk(clk),.wout(w72_30));
	PE pe72_31(.x(x31),.w(w72_30),.acc(r72_30),.res(r72_31),.clk(clk),.wout(w72_31));
	PE pe72_32(.x(x32),.w(w72_31),.acc(r72_31),.res(r72_32),.clk(clk),.wout(w72_32));
	PE pe72_33(.x(x33),.w(w72_32),.acc(r72_32),.res(r72_33),.clk(clk),.wout(w72_33));
	PE pe72_34(.x(x34),.w(w72_33),.acc(r72_33),.res(r72_34),.clk(clk),.wout(w72_34));
	PE pe72_35(.x(x35),.w(w72_34),.acc(r72_34),.res(r72_35),.clk(clk),.wout(w72_35));
	PE pe72_36(.x(x36),.w(w72_35),.acc(r72_35),.res(r72_36),.clk(clk),.wout(w72_36));
	PE pe72_37(.x(x37),.w(w72_36),.acc(r72_36),.res(r72_37),.clk(clk),.wout(w72_37));
	PE pe72_38(.x(x38),.w(w72_37),.acc(r72_37),.res(r72_38),.clk(clk),.wout(w72_38));
	PE pe72_39(.x(x39),.w(w72_38),.acc(r72_38),.res(r72_39),.clk(clk),.wout(w72_39));
	PE pe72_40(.x(x40),.w(w72_39),.acc(r72_39),.res(r72_40),.clk(clk),.wout(w72_40));
	PE pe72_41(.x(x41),.w(w72_40),.acc(r72_40),.res(r72_41),.clk(clk),.wout(w72_41));
	PE pe72_42(.x(x42),.w(w72_41),.acc(r72_41),.res(r72_42),.clk(clk),.wout(w72_42));
	PE pe72_43(.x(x43),.w(w72_42),.acc(r72_42),.res(r72_43),.clk(clk),.wout(w72_43));
	PE pe72_44(.x(x44),.w(w72_43),.acc(r72_43),.res(r72_44),.clk(clk),.wout(w72_44));
	PE pe72_45(.x(x45),.w(w72_44),.acc(r72_44),.res(r72_45),.clk(clk),.wout(w72_45));
	PE pe72_46(.x(x46),.w(w72_45),.acc(r72_45),.res(r72_46),.clk(clk),.wout(w72_46));
	PE pe72_47(.x(x47),.w(w72_46),.acc(r72_46),.res(r72_47),.clk(clk),.wout(w72_47));
	PE pe72_48(.x(x48),.w(w72_47),.acc(r72_47),.res(r72_48),.clk(clk),.wout(w72_48));
	PE pe72_49(.x(x49),.w(w72_48),.acc(r72_48),.res(r72_49),.clk(clk),.wout(w72_49));
	PE pe72_50(.x(x50),.w(w72_49),.acc(r72_49),.res(r72_50),.clk(clk),.wout(w72_50));
	PE pe72_51(.x(x51),.w(w72_50),.acc(r72_50),.res(r72_51),.clk(clk),.wout(w72_51));
	PE pe72_52(.x(x52),.w(w72_51),.acc(r72_51),.res(r72_52),.clk(clk),.wout(w72_52));
	PE pe72_53(.x(x53),.w(w72_52),.acc(r72_52),.res(r72_53),.clk(clk),.wout(w72_53));
	PE pe72_54(.x(x54),.w(w72_53),.acc(r72_53),.res(r72_54),.clk(clk),.wout(w72_54));
	PE pe72_55(.x(x55),.w(w72_54),.acc(r72_54),.res(r72_55),.clk(clk),.wout(w72_55));
	PE pe72_56(.x(x56),.w(w72_55),.acc(r72_55),.res(r72_56),.clk(clk),.wout(w72_56));
	PE pe72_57(.x(x57),.w(w72_56),.acc(r72_56),.res(r72_57),.clk(clk),.wout(w72_57));
	PE pe72_58(.x(x58),.w(w72_57),.acc(r72_57),.res(r72_58),.clk(clk),.wout(w72_58));
	PE pe72_59(.x(x59),.w(w72_58),.acc(r72_58),.res(r72_59),.clk(clk),.wout(w72_59));
	PE pe72_60(.x(x60),.w(w72_59),.acc(r72_59),.res(r72_60),.clk(clk),.wout(w72_60));
	PE pe72_61(.x(x61),.w(w72_60),.acc(r72_60),.res(r72_61),.clk(clk),.wout(w72_61));
	PE pe72_62(.x(x62),.w(w72_61),.acc(r72_61),.res(r72_62),.clk(clk),.wout(w72_62));
	PE pe72_63(.x(x63),.w(w72_62),.acc(r72_62),.res(r72_63),.clk(clk),.wout(w72_63));
	PE pe72_64(.x(x64),.w(w72_63),.acc(r72_63),.res(r72_64),.clk(clk),.wout(w72_64));
	PE pe72_65(.x(x65),.w(w72_64),.acc(r72_64),.res(r72_65),.clk(clk),.wout(w72_65));
	PE pe72_66(.x(x66),.w(w72_65),.acc(r72_65),.res(r72_66),.clk(clk),.wout(w72_66));
	PE pe72_67(.x(x67),.w(w72_66),.acc(r72_66),.res(r72_67),.clk(clk),.wout(w72_67));
	PE pe72_68(.x(x68),.w(w72_67),.acc(r72_67),.res(r72_68),.clk(clk),.wout(w72_68));
	PE pe72_69(.x(x69),.w(w72_68),.acc(r72_68),.res(r72_69),.clk(clk),.wout(w72_69));
	PE pe72_70(.x(x70),.w(w72_69),.acc(r72_69),.res(r72_70),.clk(clk),.wout(w72_70));
	PE pe72_71(.x(x71),.w(w72_70),.acc(r72_70),.res(r72_71),.clk(clk),.wout(w72_71));
	PE pe72_72(.x(x72),.w(w72_71),.acc(r72_71),.res(r72_72),.clk(clk),.wout(w72_72));
	PE pe72_73(.x(x73),.w(w72_72),.acc(r72_72),.res(r72_73),.clk(clk),.wout(w72_73));
	PE pe72_74(.x(x74),.w(w72_73),.acc(r72_73),.res(r72_74),.clk(clk),.wout(w72_74));
	PE pe72_75(.x(x75),.w(w72_74),.acc(r72_74),.res(r72_75),.clk(clk),.wout(w72_75));
	PE pe72_76(.x(x76),.w(w72_75),.acc(r72_75),.res(r72_76),.clk(clk),.wout(w72_76));
	PE pe72_77(.x(x77),.w(w72_76),.acc(r72_76),.res(r72_77),.clk(clk),.wout(w72_77));
	PE pe72_78(.x(x78),.w(w72_77),.acc(r72_77),.res(r72_78),.clk(clk),.wout(w72_78));
	PE pe72_79(.x(x79),.w(w72_78),.acc(r72_78),.res(r72_79),.clk(clk),.wout(w72_79));
	PE pe72_80(.x(x80),.w(w72_79),.acc(r72_79),.res(r72_80),.clk(clk),.wout(w72_80));
	PE pe72_81(.x(x81),.w(w72_80),.acc(r72_80),.res(r72_81),.clk(clk),.wout(w72_81));
	PE pe72_82(.x(x82),.w(w72_81),.acc(r72_81),.res(r72_82),.clk(clk),.wout(w72_82));
	PE pe72_83(.x(x83),.w(w72_82),.acc(r72_82),.res(r72_83),.clk(clk),.wout(w72_83));
	PE pe72_84(.x(x84),.w(w72_83),.acc(r72_83),.res(r72_84),.clk(clk),.wout(w72_84));
	PE pe72_85(.x(x85),.w(w72_84),.acc(r72_84),.res(r72_85),.clk(clk),.wout(w72_85));
	PE pe72_86(.x(x86),.w(w72_85),.acc(r72_85),.res(r72_86),.clk(clk),.wout(w72_86));
	PE pe72_87(.x(x87),.w(w72_86),.acc(r72_86),.res(r72_87),.clk(clk),.wout(w72_87));
	PE pe72_88(.x(x88),.w(w72_87),.acc(r72_87),.res(r72_88),.clk(clk),.wout(w72_88));
	PE pe72_89(.x(x89),.w(w72_88),.acc(r72_88),.res(r72_89),.clk(clk),.wout(w72_89));
	PE pe72_90(.x(x90),.w(w72_89),.acc(r72_89),.res(r72_90),.clk(clk),.wout(w72_90));
	PE pe72_91(.x(x91),.w(w72_90),.acc(r72_90),.res(r72_91),.clk(clk),.wout(w72_91));
	PE pe72_92(.x(x92),.w(w72_91),.acc(r72_91),.res(r72_92),.clk(clk),.wout(w72_92));
	PE pe72_93(.x(x93),.w(w72_92),.acc(r72_92),.res(r72_93),.clk(clk),.wout(w72_93));
	PE pe72_94(.x(x94),.w(w72_93),.acc(r72_93),.res(r72_94),.clk(clk),.wout(w72_94));
	PE pe72_95(.x(x95),.w(w72_94),.acc(r72_94),.res(r72_95),.clk(clk),.wout(w72_95));
	PE pe72_96(.x(x96),.w(w72_95),.acc(r72_95),.res(r72_96),.clk(clk),.wout(w72_96));
	PE pe72_97(.x(x97),.w(w72_96),.acc(r72_96),.res(r72_97),.clk(clk),.wout(w72_97));
	PE pe72_98(.x(x98),.w(w72_97),.acc(r72_97),.res(r72_98),.clk(clk),.wout(w72_98));
	PE pe72_99(.x(x99),.w(w72_98),.acc(r72_98),.res(r72_99),.clk(clk),.wout(w72_99));
	PE pe72_100(.x(x100),.w(w72_99),.acc(r72_99),.res(r72_100),.clk(clk),.wout(w72_100));
	PE pe72_101(.x(x101),.w(w72_100),.acc(r72_100),.res(r72_101),.clk(clk),.wout(w72_101));
	PE pe72_102(.x(x102),.w(w72_101),.acc(r72_101),.res(r72_102),.clk(clk),.wout(w72_102));
	PE pe72_103(.x(x103),.w(w72_102),.acc(r72_102),.res(r72_103),.clk(clk),.wout(w72_103));
	PE pe72_104(.x(x104),.w(w72_103),.acc(r72_103),.res(r72_104),.clk(clk),.wout(w72_104));
	PE pe72_105(.x(x105),.w(w72_104),.acc(r72_104),.res(r72_105),.clk(clk),.wout(w72_105));
	PE pe72_106(.x(x106),.w(w72_105),.acc(r72_105),.res(r72_106),.clk(clk),.wout(w72_106));
	PE pe72_107(.x(x107),.w(w72_106),.acc(r72_106),.res(r72_107),.clk(clk),.wout(w72_107));
	PE pe72_108(.x(x108),.w(w72_107),.acc(r72_107),.res(r72_108),.clk(clk),.wout(w72_108));
	PE pe72_109(.x(x109),.w(w72_108),.acc(r72_108),.res(r72_109),.clk(clk),.wout(w72_109));
	PE pe72_110(.x(x110),.w(w72_109),.acc(r72_109),.res(r72_110),.clk(clk),.wout(w72_110));
	PE pe72_111(.x(x111),.w(w72_110),.acc(r72_110),.res(r72_111),.clk(clk),.wout(w72_111));
	PE pe72_112(.x(x112),.w(w72_111),.acc(r72_111),.res(r72_112),.clk(clk),.wout(w72_112));
	PE pe72_113(.x(x113),.w(w72_112),.acc(r72_112),.res(r72_113),.clk(clk),.wout(w72_113));
	PE pe72_114(.x(x114),.w(w72_113),.acc(r72_113),.res(r72_114),.clk(clk),.wout(w72_114));
	PE pe72_115(.x(x115),.w(w72_114),.acc(r72_114),.res(r72_115),.clk(clk),.wout(w72_115));
	PE pe72_116(.x(x116),.w(w72_115),.acc(r72_115),.res(r72_116),.clk(clk),.wout(w72_116));
	PE pe72_117(.x(x117),.w(w72_116),.acc(r72_116),.res(r72_117),.clk(clk),.wout(w72_117));
	PE pe72_118(.x(x118),.w(w72_117),.acc(r72_117),.res(r72_118),.clk(clk),.wout(w72_118));
	PE pe72_119(.x(x119),.w(w72_118),.acc(r72_118),.res(r72_119),.clk(clk),.wout(w72_119));
	PE pe72_120(.x(x120),.w(w72_119),.acc(r72_119),.res(r72_120),.clk(clk),.wout(w72_120));
	PE pe72_121(.x(x121),.w(w72_120),.acc(r72_120),.res(r72_121),.clk(clk),.wout(w72_121));
	PE pe72_122(.x(x122),.w(w72_121),.acc(r72_121),.res(r72_122),.clk(clk),.wout(w72_122));
	PE pe72_123(.x(x123),.w(w72_122),.acc(r72_122),.res(r72_123),.clk(clk),.wout(w72_123));
	PE pe72_124(.x(x124),.w(w72_123),.acc(r72_123),.res(r72_124),.clk(clk),.wout(w72_124));
	PE pe72_125(.x(x125),.w(w72_124),.acc(r72_124),.res(r72_125),.clk(clk),.wout(w72_125));
	PE pe72_126(.x(x126),.w(w72_125),.acc(r72_125),.res(r72_126),.clk(clk),.wout(w72_126));
	PE pe72_127(.x(x127),.w(w72_126),.acc(r72_126),.res(result72),.clk(clk),.wout(weight72));

	PE pe73_0(.x(x0),.w(w73),.acc(32'h0),.res(r73_0),.clk(clk),.wout(w73_0));
	PE pe73_1(.x(x1),.w(w73_0),.acc(r73_0),.res(r73_1),.clk(clk),.wout(w73_1));
	PE pe73_2(.x(x2),.w(w73_1),.acc(r73_1),.res(r73_2),.clk(clk),.wout(w73_2));
	PE pe73_3(.x(x3),.w(w73_2),.acc(r73_2),.res(r73_3),.clk(clk),.wout(w73_3));
	PE pe73_4(.x(x4),.w(w73_3),.acc(r73_3),.res(r73_4),.clk(clk),.wout(w73_4));
	PE pe73_5(.x(x5),.w(w73_4),.acc(r73_4),.res(r73_5),.clk(clk),.wout(w73_5));
	PE pe73_6(.x(x6),.w(w73_5),.acc(r73_5),.res(r73_6),.clk(clk),.wout(w73_6));
	PE pe73_7(.x(x7),.w(w73_6),.acc(r73_6),.res(r73_7),.clk(clk),.wout(w73_7));
	PE pe73_8(.x(x8),.w(w73_7),.acc(r73_7),.res(r73_8),.clk(clk),.wout(w73_8));
	PE pe73_9(.x(x9),.w(w73_8),.acc(r73_8),.res(r73_9),.clk(clk),.wout(w73_9));
	PE pe73_10(.x(x10),.w(w73_9),.acc(r73_9),.res(r73_10),.clk(clk),.wout(w73_10));
	PE pe73_11(.x(x11),.w(w73_10),.acc(r73_10),.res(r73_11),.clk(clk),.wout(w73_11));
	PE pe73_12(.x(x12),.w(w73_11),.acc(r73_11),.res(r73_12),.clk(clk),.wout(w73_12));
	PE pe73_13(.x(x13),.w(w73_12),.acc(r73_12),.res(r73_13),.clk(clk),.wout(w73_13));
	PE pe73_14(.x(x14),.w(w73_13),.acc(r73_13),.res(r73_14),.clk(clk),.wout(w73_14));
	PE pe73_15(.x(x15),.w(w73_14),.acc(r73_14),.res(r73_15),.clk(clk),.wout(w73_15));
	PE pe73_16(.x(x16),.w(w73_15),.acc(r73_15),.res(r73_16),.clk(clk),.wout(w73_16));
	PE pe73_17(.x(x17),.w(w73_16),.acc(r73_16),.res(r73_17),.clk(clk),.wout(w73_17));
	PE pe73_18(.x(x18),.w(w73_17),.acc(r73_17),.res(r73_18),.clk(clk),.wout(w73_18));
	PE pe73_19(.x(x19),.w(w73_18),.acc(r73_18),.res(r73_19),.clk(clk),.wout(w73_19));
	PE pe73_20(.x(x20),.w(w73_19),.acc(r73_19),.res(r73_20),.clk(clk),.wout(w73_20));
	PE pe73_21(.x(x21),.w(w73_20),.acc(r73_20),.res(r73_21),.clk(clk),.wout(w73_21));
	PE pe73_22(.x(x22),.w(w73_21),.acc(r73_21),.res(r73_22),.clk(clk),.wout(w73_22));
	PE pe73_23(.x(x23),.w(w73_22),.acc(r73_22),.res(r73_23),.clk(clk),.wout(w73_23));
	PE pe73_24(.x(x24),.w(w73_23),.acc(r73_23),.res(r73_24),.clk(clk),.wout(w73_24));
	PE pe73_25(.x(x25),.w(w73_24),.acc(r73_24),.res(r73_25),.clk(clk),.wout(w73_25));
	PE pe73_26(.x(x26),.w(w73_25),.acc(r73_25),.res(r73_26),.clk(clk),.wout(w73_26));
	PE pe73_27(.x(x27),.w(w73_26),.acc(r73_26),.res(r73_27),.clk(clk),.wout(w73_27));
	PE pe73_28(.x(x28),.w(w73_27),.acc(r73_27),.res(r73_28),.clk(clk),.wout(w73_28));
	PE pe73_29(.x(x29),.w(w73_28),.acc(r73_28),.res(r73_29),.clk(clk),.wout(w73_29));
	PE pe73_30(.x(x30),.w(w73_29),.acc(r73_29),.res(r73_30),.clk(clk),.wout(w73_30));
	PE pe73_31(.x(x31),.w(w73_30),.acc(r73_30),.res(r73_31),.clk(clk),.wout(w73_31));
	PE pe73_32(.x(x32),.w(w73_31),.acc(r73_31),.res(r73_32),.clk(clk),.wout(w73_32));
	PE pe73_33(.x(x33),.w(w73_32),.acc(r73_32),.res(r73_33),.clk(clk),.wout(w73_33));
	PE pe73_34(.x(x34),.w(w73_33),.acc(r73_33),.res(r73_34),.clk(clk),.wout(w73_34));
	PE pe73_35(.x(x35),.w(w73_34),.acc(r73_34),.res(r73_35),.clk(clk),.wout(w73_35));
	PE pe73_36(.x(x36),.w(w73_35),.acc(r73_35),.res(r73_36),.clk(clk),.wout(w73_36));
	PE pe73_37(.x(x37),.w(w73_36),.acc(r73_36),.res(r73_37),.clk(clk),.wout(w73_37));
	PE pe73_38(.x(x38),.w(w73_37),.acc(r73_37),.res(r73_38),.clk(clk),.wout(w73_38));
	PE pe73_39(.x(x39),.w(w73_38),.acc(r73_38),.res(r73_39),.clk(clk),.wout(w73_39));
	PE pe73_40(.x(x40),.w(w73_39),.acc(r73_39),.res(r73_40),.clk(clk),.wout(w73_40));
	PE pe73_41(.x(x41),.w(w73_40),.acc(r73_40),.res(r73_41),.clk(clk),.wout(w73_41));
	PE pe73_42(.x(x42),.w(w73_41),.acc(r73_41),.res(r73_42),.clk(clk),.wout(w73_42));
	PE pe73_43(.x(x43),.w(w73_42),.acc(r73_42),.res(r73_43),.clk(clk),.wout(w73_43));
	PE pe73_44(.x(x44),.w(w73_43),.acc(r73_43),.res(r73_44),.clk(clk),.wout(w73_44));
	PE pe73_45(.x(x45),.w(w73_44),.acc(r73_44),.res(r73_45),.clk(clk),.wout(w73_45));
	PE pe73_46(.x(x46),.w(w73_45),.acc(r73_45),.res(r73_46),.clk(clk),.wout(w73_46));
	PE pe73_47(.x(x47),.w(w73_46),.acc(r73_46),.res(r73_47),.clk(clk),.wout(w73_47));
	PE pe73_48(.x(x48),.w(w73_47),.acc(r73_47),.res(r73_48),.clk(clk),.wout(w73_48));
	PE pe73_49(.x(x49),.w(w73_48),.acc(r73_48),.res(r73_49),.clk(clk),.wout(w73_49));
	PE pe73_50(.x(x50),.w(w73_49),.acc(r73_49),.res(r73_50),.clk(clk),.wout(w73_50));
	PE pe73_51(.x(x51),.w(w73_50),.acc(r73_50),.res(r73_51),.clk(clk),.wout(w73_51));
	PE pe73_52(.x(x52),.w(w73_51),.acc(r73_51),.res(r73_52),.clk(clk),.wout(w73_52));
	PE pe73_53(.x(x53),.w(w73_52),.acc(r73_52),.res(r73_53),.clk(clk),.wout(w73_53));
	PE pe73_54(.x(x54),.w(w73_53),.acc(r73_53),.res(r73_54),.clk(clk),.wout(w73_54));
	PE pe73_55(.x(x55),.w(w73_54),.acc(r73_54),.res(r73_55),.clk(clk),.wout(w73_55));
	PE pe73_56(.x(x56),.w(w73_55),.acc(r73_55),.res(r73_56),.clk(clk),.wout(w73_56));
	PE pe73_57(.x(x57),.w(w73_56),.acc(r73_56),.res(r73_57),.clk(clk),.wout(w73_57));
	PE pe73_58(.x(x58),.w(w73_57),.acc(r73_57),.res(r73_58),.clk(clk),.wout(w73_58));
	PE pe73_59(.x(x59),.w(w73_58),.acc(r73_58),.res(r73_59),.clk(clk),.wout(w73_59));
	PE pe73_60(.x(x60),.w(w73_59),.acc(r73_59),.res(r73_60),.clk(clk),.wout(w73_60));
	PE pe73_61(.x(x61),.w(w73_60),.acc(r73_60),.res(r73_61),.clk(clk),.wout(w73_61));
	PE pe73_62(.x(x62),.w(w73_61),.acc(r73_61),.res(r73_62),.clk(clk),.wout(w73_62));
	PE pe73_63(.x(x63),.w(w73_62),.acc(r73_62),.res(r73_63),.clk(clk),.wout(w73_63));
	PE pe73_64(.x(x64),.w(w73_63),.acc(r73_63),.res(r73_64),.clk(clk),.wout(w73_64));
	PE pe73_65(.x(x65),.w(w73_64),.acc(r73_64),.res(r73_65),.clk(clk),.wout(w73_65));
	PE pe73_66(.x(x66),.w(w73_65),.acc(r73_65),.res(r73_66),.clk(clk),.wout(w73_66));
	PE pe73_67(.x(x67),.w(w73_66),.acc(r73_66),.res(r73_67),.clk(clk),.wout(w73_67));
	PE pe73_68(.x(x68),.w(w73_67),.acc(r73_67),.res(r73_68),.clk(clk),.wout(w73_68));
	PE pe73_69(.x(x69),.w(w73_68),.acc(r73_68),.res(r73_69),.clk(clk),.wout(w73_69));
	PE pe73_70(.x(x70),.w(w73_69),.acc(r73_69),.res(r73_70),.clk(clk),.wout(w73_70));
	PE pe73_71(.x(x71),.w(w73_70),.acc(r73_70),.res(r73_71),.clk(clk),.wout(w73_71));
	PE pe73_72(.x(x72),.w(w73_71),.acc(r73_71),.res(r73_72),.clk(clk),.wout(w73_72));
	PE pe73_73(.x(x73),.w(w73_72),.acc(r73_72),.res(r73_73),.clk(clk),.wout(w73_73));
	PE pe73_74(.x(x74),.w(w73_73),.acc(r73_73),.res(r73_74),.clk(clk),.wout(w73_74));
	PE pe73_75(.x(x75),.w(w73_74),.acc(r73_74),.res(r73_75),.clk(clk),.wout(w73_75));
	PE pe73_76(.x(x76),.w(w73_75),.acc(r73_75),.res(r73_76),.clk(clk),.wout(w73_76));
	PE pe73_77(.x(x77),.w(w73_76),.acc(r73_76),.res(r73_77),.clk(clk),.wout(w73_77));
	PE pe73_78(.x(x78),.w(w73_77),.acc(r73_77),.res(r73_78),.clk(clk),.wout(w73_78));
	PE pe73_79(.x(x79),.w(w73_78),.acc(r73_78),.res(r73_79),.clk(clk),.wout(w73_79));
	PE pe73_80(.x(x80),.w(w73_79),.acc(r73_79),.res(r73_80),.clk(clk),.wout(w73_80));
	PE pe73_81(.x(x81),.w(w73_80),.acc(r73_80),.res(r73_81),.clk(clk),.wout(w73_81));
	PE pe73_82(.x(x82),.w(w73_81),.acc(r73_81),.res(r73_82),.clk(clk),.wout(w73_82));
	PE pe73_83(.x(x83),.w(w73_82),.acc(r73_82),.res(r73_83),.clk(clk),.wout(w73_83));
	PE pe73_84(.x(x84),.w(w73_83),.acc(r73_83),.res(r73_84),.clk(clk),.wout(w73_84));
	PE pe73_85(.x(x85),.w(w73_84),.acc(r73_84),.res(r73_85),.clk(clk),.wout(w73_85));
	PE pe73_86(.x(x86),.w(w73_85),.acc(r73_85),.res(r73_86),.clk(clk),.wout(w73_86));
	PE pe73_87(.x(x87),.w(w73_86),.acc(r73_86),.res(r73_87),.clk(clk),.wout(w73_87));
	PE pe73_88(.x(x88),.w(w73_87),.acc(r73_87),.res(r73_88),.clk(clk),.wout(w73_88));
	PE pe73_89(.x(x89),.w(w73_88),.acc(r73_88),.res(r73_89),.clk(clk),.wout(w73_89));
	PE pe73_90(.x(x90),.w(w73_89),.acc(r73_89),.res(r73_90),.clk(clk),.wout(w73_90));
	PE pe73_91(.x(x91),.w(w73_90),.acc(r73_90),.res(r73_91),.clk(clk),.wout(w73_91));
	PE pe73_92(.x(x92),.w(w73_91),.acc(r73_91),.res(r73_92),.clk(clk),.wout(w73_92));
	PE pe73_93(.x(x93),.w(w73_92),.acc(r73_92),.res(r73_93),.clk(clk),.wout(w73_93));
	PE pe73_94(.x(x94),.w(w73_93),.acc(r73_93),.res(r73_94),.clk(clk),.wout(w73_94));
	PE pe73_95(.x(x95),.w(w73_94),.acc(r73_94),.res(r73_95),.clk(clk),.wout(w73_95));
	PE pe73_96(.x(x96),.w(w73_95),.acc(r73_95),.res(r73_96),.clk(clk),.wout(w73_96));
	PE pe73_97(.x(x97),.w(w73_96),.acc(r73_96),.res(r73_97),.clk(clk),.wout(w73_97));
	PE pe73_98(.x(x98),.w(w73_97),.acc(r73_97),.res(r73_98),.clk(clk),.wout(w73_98));
	PE pe73_99(.x(x99),.w(w73_98),.acc(r73_98),.res(r73_99),.clk(clk),.wout(w73_99));
	PE pe73_100(.x(x100),.w(w73_99),.acc(r73_99),.res(r73_100),.clk(clk),.wout(w73_100));
	PE pe73_101(.x(x101),.w(w73_100),.acc(r73_100),.res(r73_101),.clk(clk),.wout(w73_101));
	PE pe73_102(.x(x102),.w(w73_101),.acc(r73_101),.res(r73_102),.clk(clk),.wout(w73_102));
	PE pe73_103(.x(x103),.w(w73_102),.acc(r73_102),.res(r73_103),.clk(clk),.wout(w73_103));
	PE pe73_104(.x(x104),.w(w73_103),.acc(r73_103),.res(r73_104),.clk(clk),.wout(w73_104));
	PE pe73_105(.x(x105),.w(w73_104),.acc(r73_104),.res(r73_105),.clk(clk),.wout(w73_105));
	PE pe73_106(.x(x106),.w(w73_105),.acc(r73_105),.res(r73_106),.clk(clk),.wout(w73_106));
	PE pe73_107(.x(x107),.w(w73_106),.acc(r73_106),.res(r73_107),.clk(clk),.wout(w73_107));
	PE pe73_108(.x(x108),.w(w73_107),.acc(r73_107),.res(r73_108),.clk(clk),.wout(w73_108));
	PE pe73_109(.x(x109),.w(w73_108),.acc(r73_108),.res(r73_109),.clk(clk),.wout(w73_109));
	PE pe73_110(.x(x110),.w(w73_109),.acc(r73_109),.res(r73_110),.clk(clk),.wout(w73_110));
	PE pe73_111(.x(x111),.w(w73_110),.acc(r73_110),.res(r73_111),.clk(clk),.wout(w73_111));
	PE pe73_112(.x(x112),.w(w73_111),.acc(r73_111),.res(r73_112),.clk(clk),.wout(w73_112));
	PE pe73_113(.x(x113),.w(w73_112),.acc(r73_112),.res(r73_113),.clk(clk),.wout(w73_113));
	PE pe73_114(.x(x114),.w(w73_113),.acc(r73_113),.res(r73_114),.clk(clk),.wout(w73_114));
	PE pe73_115(.x(x115),.w(w73_114),.acc(r73_114),.res(r73_115),.clk(clk),.wout(w73_115));
	PE pe73_116(.x(x116),.w(w73_115),.acc(r73_115),.res(r73_116),.clk(clk),.wout(w73_116));
	PE pe73_117(.x(x117),.w(w73_116),.acc(r73_116),.res(r73_117),.clk(clk),.wout(w73_117));
	PE pe73_118(.x(x118),.w(w73_117),.acc(r73_117),.res(r73_118),.clk(clk),.wout(w73_118));
	PE pe73_119(.x(x119),.w(w73_118),.acc(r73_118),.res(r73_119),.clk(clk),.wout(w73_119));
	PE pe73_120(.x(x120),.w(w73_119),.acc(r73_119),.res(r73_120),.clk(clk),.wout(w73_120));
	PE pe73_121(.x(x121),.w(w73_120),.acc(r73_120),.res(r73_121),.clk(clk),.wout(w73_121));
	PE pe73_122(.x(x122),.w(w73_121),.acc(r73_121),.res(r73_122),.clk(clk),.wout(w73_122));
	PE pe73_123(.x(x123),.w(w73_122),.acc(r73_122),.res(r73_123),.clk(clk),.wout(w73_123));
	PE pe73_124(.x(x124),.w(w73_123),.acc(r73_123),.res(r73_124),.clk(clk),.wout(w73_124));
	PE pe73_125(.x(x125),.w(w73_124),.acc(r73_124),.res(r73_125),.clk(clk),.wout(w73_125));
	PE pe73_126(.x(x126),.w(w73_125),.acc(r73_125),.res(r73_126),.clk(clk),.wout(w73_126));
	PE pe73_127(.x(x127),.w(w73_126),.acc(r73_126),.res(result73),.clk(clk),.wout(weight73));

	PE pe74_0(.x(x0),.w(w74),.acc(32'h0),.res(r74_0),.clk(clk),.wout(w74_0));
	PE pe74_1(.x(x1),.w(w74_0),.acc(r74_0),.res(r74_1),.clk(clk),.wout(w74_1));
	PE pe74_2(.x(x2),.w(w74_1),.acc(r74_1),.res(r74_2),.clk(clk),.wout(w74_2));
	PE pe74_3(.x(x3),.w(w74_2),.acc(r74_2),.res(r74_3),.clk(clk),.wout(w74_3));
	PE pe74_4(.x(x4),.w(w74_3),.acc(r74_3),.res(r74_4),.clk(clk),.wout(w74_4));
	PE pe74_5(.x(x5),.w(w74_4),.acc(r74_4),.res(r74_5),.clk(clk),.wout(w74_5));
	PE pe74_6(.x(x6),.w(w74_5),.acc(r74_5),.res(r74_6),.clk(clk),.wout(w74_6));
	PE pe74_7(.x(x7),.w(w74_6),.acc(r74_6),.res(r74_7),.clk(clk),.wout(w74_7));
	PE pe74_8(.x(x8),.w(w74_7),.acc(r74_7),.res(r74_8),.clk(clk),.wout(w74_8));
	PE pe74_9(.x(x9),.w(w74_8),.acc(r74_8),.res(r74_9),.clk(clk),.wout(w74_9));
	PE pe74_10(.x(x10),.w(w74_9),.acc(r74_9),.res(r74_10),.clk(clk),.wout(w74_10));
	PE pe74_11(.x(x11),.w(w74_10),.acc(r74_10),.res(r74_11),.clk(clk),.wout(w74_11));
	PE pe74_12(.x(x12),.w(w74_11),.acc(r74_11),.res(r74_12),.clk(clk),.wout(w74_12));
	PE pe74_13(.x(x13),.w(w74_12),.acc(r74_12),.res(r74_13),.clk(clk),.wout(w74_13));
	PE pe74_14(.x(x14),.w(w74_13),.acc(r74_13),.res(r74_14),.clk(clk),.wout(w74_14));
	PE pe74_15(.x(x15),.w(w74_14),.acc(r74_14),.res(r74_15),.clk(clk),.wout(w74_15));
	PE pe74_16(.x(x16),.w(w74_15),.acc(r74_15),.res(r74_16),.clk(clk),.wout(w74_16));
	PE pe74_17(.x(x17),.w(w74_16),.acc(r74_16),.res(r74_17),.clk(clk),.wout(w74_17));
	PE pe74_18(.x(x18),.w(w74_17),.acc(r74_17),.res(r74_18),.clk(clk),.wout(w74_18));
	PE pe74_19(.x(x19),.w(w74_18),.acc(r74_18),.res(r74_19),.clk(clk),.wout(w74_19));
	PE pe74_20(.x(x20),.w(w74_19),.acc(r74_19),.res(r74_20),.clk(clk),.wout(w74_20));
	PE pe74_21(.x(x21),.w(w74_20),.acc(r74_20),.res(r74_21),.clk(clk),.wout(w74_21));
	PE pe74_22(.x(x22),.w(w74_21),.acc(r74_21),.res(r74_22),.clk(clk),.wout(w74_22));
	PE pe74_23(.x(x23),.w(w74_22),.acc(r74_22),.res(r74_23),.clk(clk),.wout(w74_23));
	PE pe74_24(.x(x24),.w(w74_23),.acc(r74_23),.res(r74_24),.clk(clk),.wout(w74_24));
	PE pe74_25(.x(x25),.w(w74_24),.acc(r74_24),.res(r74_25),.clk(clk),.wout(w74_25));
	PE pe74_26(.x(x26),.w(w74_25),.acc(r74_25),.res(r74_26),.clk(clk),.wout(w74_26));
	PE pe74_27(.x(x27),.w(w74_26),.acc(r74_26),.res(r74_27),.clk(clk),.wout(w74_27));
	PE pe74_28(.x(x28),.w(w74_27),.acc(r74_27),.res(r74_28),.clk(clk),.wout(w74_28));
	PE pe74_29(.x(x29),.w(w74_28),.acc(r74_28),.res(r74_29),.clk(clk),.wout(w74_29));
	PE pe74_30(.x(x30),.w(w74_29),.acc(r74_29),.res(r74_30),.clk(clk),.wout(w74_30));
	PE pe74_31(.x(x31),.w(w74_30),.acc(r74_30),.res(r74_31),.clk(clk),.wout(w74_31));
	PE pe74_32(.x(x32),.w(w74_31),.acc(r74_31),.res(r74_32),.clk(clk),.wout(w74_32));
	PE pe74_33(.x(x33),.w(w74_32),.acc(r74_32),.res(r74_33),.clk(clk),.wout(w74_33));
	PE pe74_34(.x(x34),.w(w74_33),.acc(r74_33),.res(r74_34),.clk(clk),.wout(w74_34));
	PE pe74_35(.x(x35),.w(w74_34),.acc(r74_34),.res(r74_35),.clk(clk),.wout(w74_35));
	PE pe74_36(.x(x36),.w(w74_35),.acc(r74_35),.res(r74_36),.clk(clk),.wout(w74_36));
	PE pe74_37(.x(x37),.w(w74_36),.acc(r74_36),.res(r74_37),.clk(clk),.wout(w74_37));
	PE pe74_38(.x(x38),.w(w74_37),.acc(r74_37),.res(r74_38),.clk(clk),.wout(w74_38));
	PE pe74_39(.x(x39),.w(w74_38),.acc(r74_38),.res(r74_39),.clk(clk),.wout(w74_39));
	PE pe74_40(.x(x40),.w(w74_39),.acc(r74_39),.res(r74_40),.clk(clk),.wout(w74_40));
	PE pe74_41(.x(x41),.w(w74_40),.acc(r74_40),.res(r74_41),.clk(clk),.wout(w74_41));
	PE pe74_42(.x(x42),.w(w74_41),.acc(r74_41),.res(r74_42),.clk(clk),.wout(w74_42));
	PE pe74_43(.x(x43),.w(w74_42),.acc(r74_42),.res(r74_43),.clk(clk),.wout(w74_43));
	PE pe74_44(.x(x44),.w(w74_43),.acc(r74_43),.res(r74_44),.clk(clk),.wout(w74_44));
	PE pe74_45(.x(x45),.w(w74_44),.acc(r74_44),.res(r74_45),.clk(clk),.wout(w74_45));
	PE pe74_46(.x(x46),.w(w74_45),.acc(r74_45),.res(r74_46),.clk(clk),.wout(w74_46));
	PE pe74_47(.x(x47),.w(w74_46),.acc(r74_46),.res(r74_47),.clk(clk),.wout(w74_47));
	PE pe74_48(.x(x48),.w(w74_47),.acc(r74_47),.res(r74_48),.clk(clk),.wout(w74_48));
	PE pe74_49(.x(x49),.w(w74_48),.acc(r74_48),.res(r74_49),.clk(clk),.wout(w74_49));
	PE pe74_50(.x(x50),.w(w74_49),.acc(r74_49),.res(r74_50),.clk(clk),.wout(w74_50));
	PE pe74_51(.x(x51),.w(w74_50),.acc(r74_50),.res(r74_51),.clk(clk),.wout(w74_51));
	PE pe74_52(.x(x52),.w(w74_51),.acc(r74_51),.res(r74_52),.clk(clk),.wout(w74_52));
	PE pe74_53(.x(x53),.w(w74_52),.acc(r74_52),.res(r74_53),.clk(clk),.wout(w74_53));
	PE pe74_54(.x(x54),.w(w74_53),.acc(r74_53),.res(r74_54),.clk(clk),.wout(w74_54));
	PE pe74_55(.x(x55),.w(w74_54),.acc(r74_54),.res(r74_55),.clk(clk),.wout(w74_55));
	PE pe74_56(.x(x56),.w(w74_55),.acc(r74_55),.res(r74_56),.clk(clk),.wout(w74_56));
	PE pe74_57(.x(x57),.w(w74_56),.acc(r74_56),.res(r74_57),.clk(clk),.wout(w74_57));
	PE pe74_58(.x(x58),.w(w74_57),.acc(r74_57),.res(r74_58),.clk(clk),.wout(w74_58));
	PE pe74_59(.x(x59),.w(w74_58),.acc(r74_58),.res(r74_59),.clk(clk),.wout(w74_59));
	PE pe74_60(.x(x60),.w(w74_59),.acc(r74_59),.res(r74_60),.clk(clk),.wout(w74_60));
	PE pe74_61(.x(x61),.w(w74_60),.acc(r74_60),.res(r74_61),.clk(clk),.wout(w74_61));
	PE pe74_62(.x(x62),.w(w74_61),.acc(r74_61),.res(r74_62),.clk(clk),.wout(w74_62));
	PE pe74_63(.x(x63),.w(w74_62),.acc(r74_62),.res(r74_63),.clk(clk),.wout(w74_63));
	PE pe74_64(.x(x64),.w(w74_63),.acc(r74_63),.res(r74_64),.clk(clk),.wout(w74_64));
	PE pe74_65(.x(x65),.w(w74_64),.acc(r74_64),.res(r74_65),.clk(clk),.wout(w74_65));
	PE pe74_66(.x(x66),.w(w74_65),.acc(r74_65),.res(r74_66),.clk(clk),.wout(w74_66));
	PE pe74_67(.x(x67),.w(w74_66),.acc(r74_66),.res(r74_67),.clk(clk),.wout(w74_67));
	PE pe74_68(.x(x68),.w(w74_67),.acc(r74_67),.res(r74_68),.clk(clk),.wout(w74_68));
	PE pe74_69(.x(x69),.w(w74_68),.acc(r74_68),.res(r74_69),.clk(clk),.wout(w74_69));
	PE pe74_70(.x(x70),.w(w74_69),.acc(r74_69),.res(r74_70),.clk(clk),.wout(w74_70));
	PE pe74_71(.x(x71),.w(w74_70),.acc(r74_70),.res(r74_71),.clk(clk),.wout(w74_71));
	PE pe74_72(.x(x72),.w(w74_71),.acc(r74_71),.res(r74_72),.clk(clk),.wout(w74_72));
	PE pe74_73(.x(x73),.w(w74_72),.acc(r74_72),.res(r74_73),.clk(clk),.wout(w74_73));
	PE pe74_74(.x(x74),.w(w74_73),.acc(r74_73),.res(r74_74),.clk(clk),.wout(w74_74));
	PE pe74_75(.x(x75),.w(w74_74),.acc(r74_74),.res(r74_75),.clk(clk),.wout(w74_75));
	PE pe74_76(.x(x76),.w(w74_75),.acc(r74_75),.res(r74_76),.clk(clk),.wout(w74_76));
	PE pe74_77(.x(x77),.w(w74_76),.acc(r74_76),.res(r74_77),.clk(clk),.wout(w74_77));
	PE pe74_78(.x(x78),.w(w74_77),.acc(r74_77),.res(r74_78),.clk(clk),.wout(w74_78));
	PE pe74_79(.x(x79),.w(w74_78),.acc(r74_78),.res(r74_79),.clk(clk),.wout(w74_79));
	PE pe74_80(.x(x80),.w(w74_79),.acc(r74_79),.res(r74_80),.clk(clk),.wout(w74_80));
	PE pe74_81(.x(x81),.w(w74_80),.acc(r74_80),.res(r74_81),.clk(clk),.wout(w74_81));
	PE pe74_82(.x(x82),.w(w74_81),.acc(r74_81),.res(r74_82),.clk(clk),.wout(w74_82));
	PE pe74_83(.x(x83),.w(w74_82),.acc(r74_82),.res(r74_83),.clk(clk),.wout(w74_83));
	PE pe74_84(.x(x84),.w(w74_83),.acc(r74_83),.res(r74_84),.clk(clk),.wout(w74_84));
	PE pe74_85(.x(x85),.w(w74_84),.acc(r74_84),.res(r74_85),.clk(clk),.wout(w74_85));
	PE pe74_86(.x(x86),.w(w74_85),.acc(r74_85),.res(r74_86),.clk(clk),.wout(w74_86));
	PE pe74_87(.x(x87),.w(w74_86),.acc(r74_86),.res(r74_87),.clk(clk),.wout(w74_87));
	PE pe74_88(.x(x88),.w(w74_87),.acc(r74_87),.res(r74_88),.clk(clk),.wout(w74_88));
	PE pe74_89(.x(x89),.w(w74_88),.acc(r74_88),.res(r74_89),.clk(clk),.wout(w74_89));
	PE pe74_90(.x(x90),.w(w74_89),.acc(r74_89),.res(r74_90),.clk(clk),.wout(w74_90));
	PE pe74_91(.x(x91),.w(w74_90),.acc(r74_90),.res(r74_91),.clk(clk),.wout(w74_91));
	PE pe74_92(.x(x92),.w(w74_91),.acc(r74_91),.res(r74_92),.clk(clk),.wout(w74_92));
	PE pe74_93(.x(x93),.w(w74_92),.acc(r74_92),.res(r74_93),.clk(clk),.wout(w74_93));
	PE pe74_94(.x(x94),.w(w74_93),.acc(r74_93),.res(r74_94),.clk(clk),.wout(w74_94));
	PE pe74_95(.x(x95),.w(w74_94),.acc(r74_94),.res(r74_95),.clk(clk),.wout(w74_95));
	PE pe74_96(.x(x96),.w(w74_95),.acc(r74_95),.res(r74_96),.clk(clk),.wout(w74_96));
	PE pe74_97(.x(x97),.w(w74_96),.acc(r74_96),.res(r74_97),.clk(clk),.wout(w74_97));
	PE pe74_98(.x(x98),.w(w74_97),.acc(r74_97),.res(r74_98),.clk(clk),.wout(w74_98));
	PE pe74_99(.x(x99),.w(w74_98),.acc(r74_98),.res(r74_99),.clk(clk),.wout(w74_99));
	PE pe74_100(.x(x100),.w(w74_99),.acc(r74_99),.res(r74_100),.clk(clk),.wout(w74_100));
	PE pe74_101(.x(x101),.w(w74_100),.acc(r74_100),.res(r74_101),.clk(clk),.wout(w74_101));
	PE pe74_102(.x(x102),.w(w74_101),.acc(r74_101),.res(r74_102),.clk(clk),.wout(w74_102));
	PE pe74_103(.x(x103),.w(w74_102),.acc(r74_102),.res(r74_103),.clk(clk),.wout(w74_103));
	PE pe74_104(.x(x104),.w(w74_103),.acc(r74_103),.res(r74_104),.clk(clk),.wout(w74_104));
	PE pe74_105(.x(x105),.w(w74_104),.acc(r74_104),.res(r74_105),.clk(clk),.wout(w74_105));
	PE pe74_106(.x(x106),.w(w74_105),.acc(r74_105),.res(r74_106),.clk(clk),.wout(w74_106));
	PE pe74_107(.x(x107),.w(w74_106),.acc(r74_106),.res(r74_107),.clk(clk),.wout(w74_107));
	PE pe74_108(.x(x108),.w(w74_107),.acc(r74_107),.res(r74_108),.clk(clk),.wout(w74_108));
	PE pe74_109(.x(x109),.w(w74_108),.acc(r74_108),.res(r74_109),.clk(clk),.wout(w74_109));
	PE pe74_110(.x(x110),.w(w74_109),.acc(r74_109),.res(r74_110),.clk(clk),.wout(w74_110));
	PE pe74_111(.x(x111),.w(w74_110),.acc(r74_110),.res(r74_111),.clk(clk),.wout(w74_111));
	PE pe74_112(.x(x112),.w(w74_111),.acc(r74_111),.res(r74_112),.clk(clk),.wout(w74_112));
	PE pe74_113(.x(x113),.w(w74_112),.acc(r74_112),.res(r74_113),.clk(clk),.wout(w74_113));
	PE pe74_114(.x(x114),.w(w74_113),.acc(r74_113),.res(r74_114),.clk(clk),.wout(w74_114));
	PE pe74_115(.x(x115),.w(w74_114),.acc(r74_114),.res(r74_115),.clk(clk),.wout(w74_115));
	PE pe74_116(.x(x116),.w(w74_115),.acc(r74_115),.res(r74_116),.clk(clk),.wout(w74_116));
	PE pe74_117(.x(x117),.w(w74_116),.acc(r74_116),.res(r74_117),.clk(clk),.wout(w74_117));
	PE pe74_118(.x(x118),.w(w74_117),.acc(r74_117),.res(r74_118),.clk(clk),.wout(w74_118));
	PE pe74_119(.x(x119),.w(w74_118),.acc(r74_118),.res(r74_119),.clk(clk),.wout(w74_119));
	PE pe74_120(.x(x120),.w(w74_119),.acc(r74_119),.res(r74_120),.clk(clk),.wout(w74_120));
	PE pe74_121(.x(x121),.w(w74_120),.acc(r74_120),.res(r74_121),.clk(clk),.wout(w74_121));
	PE pe74_122(.x(x122),.w(w74_121),.acc(r74_121),.res(r74_122),.clk(clk),.wout(w74_122));
	PE pe74_123(.x(x123),.w(w74_122),.acc(r74_122),.res(r74_123),.clk(clk),.wout(w74_123));
	PE pe74_124(.x(x124),.w(w74_123),.acc(r74_123),.res(r74_124),.clk(clk),.wout(w74_124));
	PE pe74_125(.x(x125),.w(w74_124),.acc(r74_124),.res(r74_125),.clk(clk),.wout(w74_125));
	PE pe74_126(.x(x126),.w(w74_125),.acc(r74_125),.res(r74_126),.clk(clk),.wout(w74_126));
	PE pe74_127(.x(x127),.w(w74_126),.acc(r74_126),.res(result74),.clk(clk),.wout(weight74));

	PE pe75_0(.x(x0),.w(w75),.acc(32'h0),.res(r75_0),.clk(clk),.wout(w75_0));
	PE pe75_1(.x(x1),.w(w75_0),.acc(r75_0),.res(r75_1),.clk(clk),.wout(w75_1));
	PE pe75_2(.x(x2),.w(w75_1),.acc(r75_1),.res(r75_2),.clk(clk),.wout(w75_2));
	PE pe75_3(.x(x3),.w(w75_2),.acc(r75_2),.res(r75_3),.clk(clk),.wout(w75_3));
	PE pe75_4(.x(x4),.w(w75_3),.acc(r75_3),.res(r75_4),.clk(clk),.wout(w75_4));
	PE pe75_5(.x(x5),.w(w75_4),.acc(r75_4),.res(r75_5),.clk(clk),.wout(w75_5));
	PE pe75_6(.x(x6),.w(w75_5),.acc(r75_5),.res(r75_6),.clk(clk),.wout(w75_6));
	PE pe75_7(.x(x7),.w(w75_6),.acc(r75_6),.res(r75_7),.clk(clk),.wout(w75_7));
	PE pe75_8(.x(x8),.w(w75_7),.acc(r75_7),.res(r75_8),.clk(clk),.wout(w75_8));
	PE pe75_9(.x(x9),.w(w75_8),.acc(r75_8),.res(r75_9),.clk(clk),.wout(w75_9));
	PE pe75_10(.x(x10),.w(w75_9),.acc(r75_9),.res(r75_10),.clk(clk),.wout(w75_10));
	PE pe75_11(.x(x11),.w(w75_10),.acc(r75_10),.res(r75_11),.clk(clk),.wout(w75_11));
	PE pe75_12(.x(x12),.w(w75_11),.acc(r75_11),.res(r75_12),.clk(clk),.wout(w75_12));
	PE pe75_13(.x(x13),.w(w75_12),.acc(r75_12),.res(r75_13),.clk(clk),.wout(w75_13));
	PE pe75_14(.x(x14),.w(w75_13),.acc(r75_13),.res(r75_14),.clk(clk),.wout(w75_14));
	PE pe75_15(.x(x15),.w(w75_14),.acc(r75_14),.res(r75_15),.clk(clk),.wout(w75_15));
	PE pe75_16(.x(x16),.w(w75_15),.acc(r75_15),.res(r75_16),.clk(clk),.wout(w75_16));
	PE pe75_17(.x(x17),.w(w75_16),.acc(r75_16),.res(r75_17),.clk(clk),.wout(w75_17));
	PE pe75_18(.x(x18),.w(w75_17),.acc(r75_17),.res(r75_18),.clk(clk),.wout(w75_18));
	PE pe75_19(.x(x19),.w(w75_18),.acc(r75_18),.res(r75_19),.clk(clk),.wout(w75_19));
	PE pe75_20(.x(x20),.w(w75_19),.acc(r75_19),.res(r75_20),.clk(clk),.wout(w75_20));
	PE pe75_21(.x(x21),.w(w75_20),.acc(r75_20),.res(r75_21),.clk(clk),.wout(w75_21));
	PE pe75_22(.x(x22),.w(w75_21),.acc(r75_21),.res(r75_22),.clk(clk),.wout(w75_22));
	PE pe75_23(.x(x23),.w(w75_22),.acc(r75_22),.res(r75_23),.clk(clk),.wout(w75_23));
	PE pe75_24(.x(x24),.w(w75_23),.acc(r75_23),.res(r75_24),.clk(clk),.wout(w75_24));
	PE pe75_25(.x(x25),.w(w75_24),.acc(r75_24),.res(r75_25),.clk(clk),.wout(w75_25));
	PE pe75_26(.x(x26),.w(w75_25),.acc(r75_25),.res(r75_26),.clk(clk),.wout(w75_26));
	PE pe75_27(.x(x27),.w(w75_26),.acc(r75_26),.res(r75_27),.clk(clk),.wout(w75_27));
	PE pe75_28(.x(x28),.w(w75_27),.acc(r75_27),.res(r75_28),.clk(clk),.wout(w75_28));
	PE pe75_29(.x(x29),.w(w75_28),.acc(r75_28),.res(r75_29),.clk(clk),.wout(w75_29));
	PE pe75_30(.x(x30),.w(w75_29),.acc(r75_29),.res(r75_30),.clk(clk),.wout(w75_30));
	PE pe75_31(.x(x31),.w(w75_30),.acc(r75_30),.res(r75_31),.clk(clk),.wout(w75_31));
	PE pe75_32(.x(x32),.w(w75_31),.acc(r75_31),.res(r75_32),.clk(clk),.wout(w75_32));
	PE pe75_33(.x(x33),.w(w75_32),.acc(r75_32),.res(r75_33),.clk(clk),.wout(w75_33));
	PE pe75_34(.x(x34),.w(w75_33),.acc(r75_33),.res(r75_34),.clk(clk),.wout(w75_34));
	PE pe75_35(.x(x35),.w(w75_34),.acc(r75_34),.res(r75_35),.clk(clk),.wout(w75_35));
	PE pe75_36(.x(x36),.w(w75_35),.acc(r75_35),.res(r75_36),.clk(clk),.wout(w75_36));
	PE pe75_37(.x(x37),.w(w75_36),.acc(r75_36),.res(r75_37),.clk(clk),.wout(w75_37));
	PE pe75_38(.x(x38),.w(w75_37),.acc(r75_37),.res(r75_38),.clk(clk),.wout(w75_38));
	PE pe75_39(.x(x39),.w(w75_38),.acc(r75_38),.res(r75_39),.clk(clk),.wout(w75_39));
	PE pe75_40(.x(x40),.w(w75_39),.acc(r75_39),.res(r75_40),.clk(clk),.wout(w75_40));
	PE pe75_41(.x(x41),.w(w75_40),.acc(r75_40),.res(r75_41),.clk(clk),.wout(w75_41));
	PE pe75_42(.x(x42),.w(w75_41),.acc(r75_41),.res(r75_42),.clk(clk),.wout(w75_42));
	PE pe75_43(.x(x43),.w(w75_42),.acc(r75_42),.res(r75_43),.clk(clk),.wout(w75_43));
	PE pe75_44(.x(x44),.w(w75_43),.acc(r75_43),.res(r75_44),.clk(clk),.wout(w75_44));
	PE pe75_45(.x(x45),.w(w75_44),.acc(r75_44),.res(r75_45),.clk(clk),.wout(w75_45));
	PE pe75_46(.x(x46),.w(w75_45),.acc(r75_45),.res(r75_46),.clk(clk),.wout(w75_46));
	PE pe75_47(.x(x47),.w(w75_46),.acc(r75_46),.res(r75_47),.clk(clk),.wout(w75_47));
	PE pe75_48(.x(x48),.w(w75_47),.acc(r75_47),.res(r75_48),.clk(clk),.wout(w75_48));
	PE pe75_49(.x(x49),.w(w75_48),.acc(r75_48),.res(r75_49),.clk(clk),.wout(w75_49));
	PE pe75_50(.x(x50),.w(w75_49),.acc(r75_49),.res(r75_50),.clk(clk),.wout(w75_50));
	PE pe75_51(.x(x51),.w(w75_50),.acc(r75_50),.res(r75_51),.clk(clk),.wout(w75_51));
	PE pe75_52(.x(x52),.w(w75_51),.acc(r75_51),.res(r75_52),.clk(clk),.wout(w75_52));
	PE pe75_53(.x(x53),.w(w75_52),.acc(r75_52),.res(r75_53),.clk(clk),.wout(w75_53));
	PE pe75_54(.x(x54),.w(w75_53),.acc(r75_53),.res(r75_54),.clk(clk),.wout(w75_54));
	PE pe75_55(.x(x55),.w(w75_54),.acc(r75_54),.res(r75_55),.clk(clk),.wout(w75_55));
	PE pe75_56(.x(x56),.w(w75_55),.acc(r75_55),.res(r75_56),.clk(clk),.wout(w75_56));
	PE pe75_57(.x(x57),.w(w75_56),.acc(r75_56),.res(r75_57),.clk(clk),.wout(w75_57));
	PE pe75_58(.x(x58),.w(w75_57),.acc(r75_57),.res(r75_58),.clk(clk),.wout(w75_58));
	PE pe75_59(.x(x59),.w(w75_58),.acc(r75_58),.res(r75_59),.clk(clk),.wout(w75_59));
	PE pe75_60(.x(x60),.w(w75_59),.acc(r75_59),.res(r75_60),.clk(clk),.wout(w75_60));
	PE pe75_61(.x(x61),.w(w75_60),.acc(r75_60),.res(r75_61),.clk(clk),.wout(w75_61));
	PE pe75_62(.x(x62),.w(w75_61),.acc(r75_61),.res(r75_62),.clk(clk),.wout(w75_62));
	PE pe75_63(.x(x63),.w(w75_62),.acc(r75_62),.res(r75_63),.clk(clk),.wout(w75_63));
	PE pe75_64(.x(x64),.w(w75_63),.acc(r75_63),.res(r75_64),.clk(clk),.wout(w75_64));
	PE pe75_65(.x(x65),.w(w75_64),.acc(r75_64),.res(r75_65),.clk(clk),.wout(w75_65));
	PE pe75_66(.x(x66),.w(w75_65),.acc(r75_65),.res(r75_66),.clk(clk),.wout(w75_66));
	PE pe75_67(.x(x67),.w(w75_66),.acc(r75_66),.res(r75_67),.clk(clk),.wout(w75_67));
	PE pe75_68(.x(x68),.w(w75_67),.acc(r75_67),.res(r75_68),.clk(clk),.wout(w75_68));
	PE pe75_69(.x(x69),.w(w75_68),.acc(r75_68),.res(r75_69),.clk(clk),.wout(w75_69));
	PE pe75_70(.x(x70),.w(w75_69),.acc(r75_69),.res(r75_70),.clk(clk),.wout(w75_70));
	PE pe75_71(.x(x71),.w(w75_70),.acc(r75_70),.res(r75_71),.clk(clk),.wout(w75_71));
	PE pe75_72(.x(x72),.w(w75_71),.acc(r75_71),.res(r75_72),.clk(clk),.wout(w75_72));
	PE pe75_73(.x(x73),.w(w75_72),.acc(r75_72),.res(r75_73),.clk(clk),.wout(w75_73));
	PE pe75_74(.x(x74),.w(w75_73),.acc(r75_73),.res(r75_74),.clk(clk),.wout(w75_74));
	PE pe75_75(.x(x75),.w(w75_74),.acc(r75_74),.res(r75_75),.clk(clk),.wout(w75_75));
	PE pe75_76(.x(x76),.w(w75_75),.acc(r75_75),.res(r75_76),.clk(clk),.wout(w75_76));
	PE pe75_77(.x(x77),.w(w75_76),.acc(r75_76),.res(r75_77),.clk(clk),.wout(w75_77));
	PE pe75_78(.x(x78),.w(w75_77),.acc(r75_77),.res(r75_78),.clk(clk),.wout(w75_78));
	PE pe75_79(.x(x79),.w(w75_78),.acc(r75_78),.res(r75_79),.clk(clk),.wout(w75_79));
	PE pe75_80(.x(x80),.w(w75_79),.acc(r75_79),.res(r75_80),.clk(clk),.wout(w75_80));
	PE pe75_81(.x(x81),.w(w75_80),.acc(r75_80),.res(r75_81),.clk(clk),.wout(w75_81));
	PE pe75_82(.x(x82),.w(w75_81),.acc(r75_81),.res(r75_82),.clk(clk),.wout(w75_82));
	PE pe75_83(.x(x83),.w(w75_82),.acc(r75_82),.res(r75_83),.clk(clk),.wout(w75_83));
	PE pe75_84(.x(x84),.w(w75_83),.acc(r75_83),.res(r75_84),.clk(clk),.wout(w75_84));
	PE pe75_85(.x(x85),.w(w75_84),.acc(r75_84),.res(r75_85),.clk(clk),.wout(w75_85));
	PE pe75_86(.x(x86),.w(w75_85),.acc(r75_85),.res(r75_86),.clk(clk),.wout(w75_86));
	PE pe75_87(.x(x87),.w(w75_86),.acc(r75_86),.res(r75_87),.clk(clk),.wout(w75_87));
	PE pe75_88(.x(x88),.w(w75_87),.acc(r75_87),.res(r75_88),.clk(clk),.wout(w75_88));
	PE pe75_89(.x(x89),.w(w75_88),.acc(r75_88),.res(r75_89),.clk(clk),.wout(w75_89));
	PE pe75_90(.x(x90),.w(w75_89),.acc(r75_89),.res(r75_90),.clk(clk),.wout(w75_90));
	PE pe75_91(.x(x91),.w(w75_90),.acc(r75_90),.res(r75_91),.clk(clk),.wout(w75_91));
	PE pe75_92(.x(x92),.w(w75_91),.acc(r75_91),.res(r75_92),.clk(clk),.wout(w75_92));
	PE pe75_93(.x(x93),.w(w75_92),.acc(r75_92),.res(r75_93),.clk(clk),.wout(w75_93));
	PE pe75_94(.x(x94),.w(w75_93),.acc(r75_93),.res(r75_94),.clk(clk),.wout(w75_94));
	PE pe75_95(.x(x95),.w(w75_94),.acc(r75_94),.res(r75_95),.clk(clk),.wout(w75_95));
	PE pe75_96(.x(x96),.w(w75_95),.acc(r75_95),.res(r75_96),.clk(clk),.wout(w75_96));
	PE pe75_97(.x(x97),.w(w75_96),.acc(r75_96),.res(r75_97),.clk(clk),.wout(w75_97));
	PE pe75_98(.x(x98),.w(w75_97),.acc(r75_97),.res(r75_98),.clk(clk),.wout(w75_98));
	PE pe75_99(.x(x99),.w(w75_98),.acc(r75_98),.res(r75_99),.clk(clk),.wout(w75_99));
	PE pe75_100(.x(x100),.w(w75_99),.acc(r75_99),.res(r75_100),.clk(clk),.wout(w75_100));
	PE pe75_101(.x(x101),.w(w75_100),.acc(r75_100),.res(r75_101),.clk(clk),.wout(w75_101));
	PE pe75_102(.x(x102),.w(w75_101),.acc(r75_101),.res(r75_102),.clk(clk),.wout(w75_102));
	PE pe75_103(.x(x103),.w(w75_102),.acc(r75_102),.res(r75_103),.clk(clk),.wout(w75_103));
	PE pe75_104(.x(x104),.w(w75_103),.acc(r75_103),.res(r75_104),.clk(clk),.wout(w75_104));
	PE pe75_105(.x(x105),.w(w75_104),.acc(r75_104),.res(r75_105),.clk(clk),.wout(w75_105));
	PE pe75_106(.x(x106),.w(w75_105),.acc(r75_105),.res(r75_106),.clk(clk),.wout(w75_106));
	PE pe75_107(.x(x107),.w(w75_106),.acc(r75_106),.res(r75_107),.clk(clk),.wout(w75_107));
	PE pe75_108(.x(x108),.w(w75_107),.acc(r75_107),.res(r75_108),.clk(clk),.wout(w75_108));
	PE pe75_109(.x(x109),.w(w75_108),.acc(r75_108),.res(r75_109),.clk(clk),.wout(w75_109));
	PE pe75_110(.x(x110),.w(w75_109),.acc(r75_109),.res(r75_110),.clk(clk),.wout(w75_110));
	PE pe75_111(.x(x111),.w(w75_110),.acc(r75_110),.res(r75_111),.clk(clk),.wout(w75_111));
	PE pe75_112(.x(x112),.w(w75_111),.acc(r75_111),.res(r75_112),.clk(clk),.wout(w75_112));
	PE pe75_113(.x(x113),.w(w75_112),.acc(r75_112),.res(r75_113),.clk(clk),.wout(w75_113));
	PE pe75_114(.x(x114),.w(w75_113),.acc(r75_113),.res(r75_114),.clk(clk),.wout(w75_114));
	PE pe75_115(.x(x115),.w(w75_114),.acc(r75_114),.res(r75_115),.clk(clk),.wout(w75_115));
	PE pe75_116(.x(x116),.w(w75_115),.acc(r75_115),.res(r75_116),.clk(clk),.wout(w75_116));
	PE pe75_117(.x(x117),.w(w75_116),.acc(r75_116),.res(r75_117),.clk(clk),.wout(w75_117));
	PE pe75_118(.x(x118),.w(w75_117),.acc(r75_117),.res(r75_118),.clk(clk),.wout(w75_118));
	PE pe75_119(.x(x119),.w(w75_118),.acc(r75_118),.res(r75_119),.clk(clk),.wout(w75_119));
	PE pe75_120(.x(x120),.w(w75_119),.acc(r75_119),.res(r75_120),.clk(clk),.wout(w75_120));
	PE pe75_121(.x(x121),.w(w75_120),.acc(r75_120),.res(r75_121),.clk(clk),.wout(w75_121));
	PE pe75_122(.x(x122),.w(w75_121),.acc(r75_121),.res(r75_122),.clk(clk),.wout(w75_122));
	PE pe75_123(.x(x123),.w(w75_122),.acc(r75_122),.res(r75_123),.clk(clk),.wout(w75_123));
	PE pe75_124(.x(x124),.w(w75_123),.acc(r75_123),.res(r75_124),.clk(clk),.wout(w75_124));
	PE pe75_125(.x(x125),.w(w75_124),.acc(r75_124),.res(r75_125),.clk(clk),.wout(w75_125));
	PE pe75_126(.x(x126),.w(w75_125),.acc(r75_125),.res(r75_126),.clk(clk),.wout(w75_126));
	PE pe75_127(.x(x127),.w(w75_126),.acc(r75_126),.res(result75),.clk(clk),.wout(weight75));

	PE pe76_0(.x(x0),.w(w76),.acc(32'h0),.res(r76_0),.clk(clk),.wout(w76_0));
	PE pe76_1(.x(x1),.w(w76_0),.acc(r76_0),.res(r76_1),.clk(clk),.wout(w76_1));
	PE pe76_2(.x(x2),.w(w76_1),.acc(r76_1),.res(r76_2),.clk(clk),.wout(w76_2));
	PE pe76_3(.x(x3),.w(w76_2),.acc(r76_2),.res(r76_3),.clk(clk),.wout(w76_3));
	PE pe76_4(.x(x4),.w(w76_3),.acc(r76_3),.res(r76_4),.clk(clk),.wout(w76_4));
	PE pe76_5(.x(x5),.w(w76_4),.acc(r76_4),.res(r76_5),.clk(clk),.wout(w76_5));
	PE pe76_6(.x(x6),.w(w76_5),.acc(r76_5),.res(r76_6),.clk(clk),.wout(w76_6));
	PE pe76_7(.x(x7),.w(w76_6),.acc(r76_6),.res(r76_7),.clk(clk),.wout(w76_7));
	PE pe76_8(.x(x8),.w(w76_7),.acc(r76_7),.res(r76_8),.clk(clk),.wout(w76_8));
	PE pe76_9(.x(x9),.w(w76_8),.acc(r76_8),.res(r76_9),.clk(clk),.wout(w76_9));
	PE pe76_10(.x(x10),.w(w76_9),.acc(r76_9),.res(r76_10),.clk(clk),.wout(w76_10));
	PE pe76_11(.x(x11),.w(w76_10),.acc(r76_10),.res(r76_11),.clk(clk),.wout(w76_11));
	PE pe76_12(.x(x12),.w(w76_11),.acc(r76_11),.res(r76_12),.clk(clk),.wout(w76_12));
	PE pe76_13(.x(x13),.w(w76_12),.acc(r76_12),.res(r76_13),.clk(clk),.wout(w76_13));
	PE pe76_14(.x(x14),.w(w76_13),.acc(r76_13),.res(r76_14),.clk(clk),.wout(w76_14));
	PE pe76_15(.x(x15),.w(w76_14),.acc(r76_14),.res(r76_15),.clk(clk),.wout(w76_15));
	PE pe76_16(.x(x16),.w(w76_15),.acc(r76_15),.res(r76_16),.clk(clk),.wout(w76_16));
	PE pe76_17(.x(x17),.w(w76_16),.acc(r76_16),.res(r76_17),.clk(clk),.wout(w76_17));
	PE pe76_18(.x(x18),.w(w76_17),.acc(r76_17),.res(r76_18),.clk(clk),.wout(w76_18));
	PE pe76_19(.x(x19),.w(w76_18),.acc(r76_18),.res(r76_19),.clk(clk),.wout(w76_19));
	PE pe76_20(.x(x20),.w(w76_19),.acc(r76_19),.res(r76_20),.clk(clk),.wout(w76_20));
	PE pe76_21(.x(x21),.w(w76_20),.acc(r76_20),.res(r76_21),.clk(clk),.wout(w76_21));
	PE pe76_22(.x(x22),.w(w76_21),.acc(r76_21),.res(r76_22),.clk(clk),.wout(w76_22));
	PE pe76_23(.x(x23),.w(w76_22),.acc(r76_22),.res(r76_23),.clk(clk),.wout(w76_23));
	PE pe76_24(.x(x24),.w(w76_23),.acc(r76_23),.res(r76_24),.clk(clk),.wout(w76_24));
	PE pe76_25(.x(x25),.w(w76_24),.acc(r76_24),.res(r76_25),.clk(clk),.wout(w76_25));
	PE pe76_26(.x(x26),.w(w76_25),.acc(r76_25),.res(r76_26),.clk(clk),.wout(w76_26));
	PE pe76_27(.x(x27),.w(w76_26),.acc(r76_26),.res(r76_27),.clk(clk),.wout(w76_27));
	PE pe76_28(.x(x28),.w(w76_27),.acc(r76_27),.res(r76_28),.clk(clk),.wout(w76_28));
	PE pe76_29(.x(x29),.w(w76_28),.acc(r76_28),.res(r76_29),.clk(clk),.wout(w76_29));
	PE pe76_30(.x(x30),.w(w76_29),.acc(r76_29),.res(r76_30),.clk(clk),.wout(w76_30));
	PE pe76_31(.x(x31),.w(w76_30),.acc(r76_30),.res(r76_31),.clk(clk),.wout(w76_31));
	PE pe76_32(.x(x32),.w(w76_31),.acc(r76_31),.res(r76_32),.clk(clk),.wout(w76_32));
	PE pe76_33(.x(x33),.w(w76_32),.acc(r76_32),.res(r76_33),.clk(clk),.wout(w76_33));
	PE pe76_34(.x(x34),.w(w76_33),.acc(r76_33),.res(r76_34),.clk(clk),.wout(w76_34));
	PE pe76_35(.x(x35),.w(w76_34),.acc(r76_34),.res(r76_35),.clk(clk),.wout(w76_35));
	PE pe76_36(.x(x36),.w(w76_35),.acc(r76_35),.res(r76_36),.clk(clk),.wout(w76_36));
	PE pe76_37(.x(x37),.w(w76_36),.acc(r76_36),.res(r76_37),.clk(clk),.wout(w76_37));
	PE pe76_38(.x(x38),.w(w76_37),.acc(r76_37),.res(r76_38),.clk(clk),.wout(w76_38));
	PE pe76_39(.x(x39),.w(w76_38),.acc(r76_38),.res(r76_39),.clk(clk),.wout(w76_39));
	PE pe76_40(.x(x40),.w(w76_39),.acc(r76_39),.res(r76_40),.clk(clk),.wout(w76_40));
	PE pe76_41(.x(x41),.w(w76_40),.acc(r76_40),.res(r76_41),.clk(clk),.wout(w76_41));
	PE pe76_42(.x(x42),.w(w76_41),.acc(r76_41),.res(r76_42),.clk(clk),.wout(w76_42));
	PE pe76_43(.x(x43),.w(w76_42),.acc(r76_42),.res(r76_43),.clk(clk),.wout(w76_43));
	PE pe76_44(.x(x44),.w(w76_43),.acc(r76_43),.res(r76_44),.clk(clk),.wout(w76_44));
	PE pe76_45(.x(x45),.w(w76_44),.acc(r76_44),.res(r76_45),.clk(clk),.wout(w76_45));
	PE pe76_46(.x(x46),.w(w76_45),.acc(r76_45),.res(r76_46),.clk(clk),.wout(w76_46));
	PE pe76_47(.x(x47),.w(w76_46),.acc(r76_46),.res(r76_47),.clk(clk),.wout(w76_47));
	PE pe76_48(.x(x48),.w(w76_47),.acc(r76_47),.res(r76_48),.clk(clk),.wout(w76_48));
	PE pe76_49(.x(x49),.w(w76_48),.acc(r76_48),.res(r76_49),.clk(clk),.wout(w76_49));
	PE pe76_50(.x(x50),.w(w76_49),.acc(r76_49),.res(r76_50),.clk(clk),.wout(w76_50));
	PE pe76_51(.x(x51),.w(w76_50),.acc(r76_50),.res(r76_51),.clk(clk),.wout(w76_51));
	PE pe76_52(.x(x52),.w(w76_51),.acc(r76_51),.res(r76_52),.clk(clk),.wout(w76_52));
	PE pe76_53(.x(x53),.w(w76_52),.acc(r76_52),.res(r76_53),.clk(clk),.wout(w76_53));
	PE pe76_54(.x(x54),.w(w76_53),.acc(r76_53),.res(r76_54),.clk(clk),.wout(w76_54));
	PE pe76_55(.x(x55),.w(w76_54),.acc(r76_54),.res(r76_55),.clk(clk),.wout(w76_55));
	PE pe76_56(.x(x56),.w(w76_55),.acc(r76_55),.res(r76_56),.clk(clk),.wout(w76_56));
	PE pe76_57(.x(x57),.w(w76_56),.acc(r76_56),.res(r76_57),.clk(clk),.wout(w76_57));
	PE pe76_58(.x(x58),.w(w76_57),.acc(r76_57),.res(r76_58),.clk(clk),.wout(w76_58));
	PE pe76_59(.x(x59),.w(w76_58),.acc(r76_58),.res(r76_59),.clk(clk),.wout(w76_59));
	PE pe76_60(.x(x60),.w(w76_59),.acc(r76_59),.res(r76_60),.clk(clk),.wout(w76_60));
	PE pe76_61(.x(x61),.w(w76_60),.acc(r76_60),.res(r76_61),.clk(clk),.wout(w76_61));
	PE pe76_62(.x(x62),.w(w76_61),.acc(r76_61),.res(r76_62),.clk(clk),.wout(w76_62));
	PE pe76_63(.x(x63),.w(w76_62),.acc(r76_62),.res(r76_63),.clk(clk),.wout(w76_63));
	PE pe76_64(.x(x64),.w(w76_63),.acc(r76_63),.res(r76_64),.clk(clk),.wout(w76_64));
	PE pe76_65(.x(x65),.w(w76_64),.acc(r76_64),.res(r76_65),.clk(clk),.wout(w76_65));
	PE pe76_66(.x(x66),.w(w76_65),.acc(r76_65),.res(r76_66),.clk(clk),.wout(w76_66));
	PE pe76_67(.x(x67),.w(w76_66),.acc(r76_66),.res(r76_67),.clk(clk),.wout(w76_67));
	PE pe76_68(.x(x68),.w(w76_67),.acc(r76_67),.res(r76_68),.clk(clk),.wout(w76_68));
	PE pe76_69(.x(x69),.w(w76_68),.acc(r76_68),.res(r76_69),.clk(clk),.wout(w76_69));
	PE pe76_70(.x(x70),.w(w76_69),.acc(r76_69),.res(r76_70),.clk(clk),.wout(w76_70));
	PE pe76_71(.x(x71),.w(w76_70),.acc(r76_70),.res(r76_71),.clk(clk),.wout(w76_71));
	PE pe76_72(.x(x72),.w(w76_71),.acc(r76_71),.res(r76_72),.clk(clk),.wout(w76_72));
	PE pe76_73(.x(x73),.w(w76_72),.acc(r76_72),.res(r76_73),.clk(clk),.wout(w76_73));
	PE pe76_74(.x(x74),.w(w76_73),.acc(r76_73),.res(r76_74),.clk(clk),.wout(w76_74));
	PE pe76_75(.x(x75),.w(w76_74),.acc(r76_74),.res(r76_75),.clk(clk),.wout(w76_75));
	PE pe76_76(.x(x76),.w(w76_75),.acc(r76_75),.res(r76_76),.clk(clk),.wout(w76_76));
	PE pe76_77(.x(x77),.w(w76_76),.acc(r76_76),.res(r76_77),.clk(clk),.wout(w76_77));
	PE pe76_78(.x(x78),.w(w76_77),.acc(r76_77),.res(r76_78),.clk(clk),.wout(w76_78));
	PE pe76_79(.x(x79),.w(w76_78),.acc(r76_78),.res(r76_79),.clk(clk),.wout(w76_79));
	PE pe76_80(.x(x80),.w(w76_79),.acc(r76_79),.res(r76_80),.clk(clk),.wout(w76_80));
	PE pe76_81(.x(x81),.w(w76_80),.acc(r76_80),.res(r76_81),.clk(clk),.wout(w76_81));
	PE pe76_82(.x(x82),.w(w76_81),.acc(r76_81),.res(r76_82),.clk(clk),.wout(w76_82));
	PE pe76_83(.x(x83),.w(w76_82),.acc(r76_82),.res(r76_83),.clk(clk),.wout(w76_83));
	PE pe76_84(.x(x84),.w(w76_83),.acc(r76_83),.res(r76_84),.clk(clk),.wout(w76_84));
	PE pe76_85(.x(x85),.w(w76_84),.acc(r76_84),.res(r76_85),.clk(clk),.wout(w76_85));
	PE pe76_86(.x(x86),.w(w76_85),.acc(r76_85),.res(r76_86),.clk(clk),.wout(w76_86));
	PE pe76_87(.x(x87),.w(w76_86),.acc(r76_86),.res(r76_87),.clk(clk),.wout(w76_87));
	PE pe76_88(.x(x88),.w(w76_87),.acc(r76_87),.res(r76_88),.clk(clk),.wout(w76_88));
	PE pe76_89(.x(x89),.w(w76_88),.acc(r76_88),.res(r76_89),.clk(clk),.wout(w76_89));
	PE pe76_90(.x(x90),.w(w76_89),.acc(r76_89),.res(r76_90),.clk(clk),.wout(w76_90));
	PE pe76_91(.x(x91),.w(w76_90),.acc(r76_90),.res(r76_91),.clk(clk),.wout(w76_91));
	PE pe76_92(.x(x92),.w(w76_91),.acc(r76_91),.res(r76_92),.clk(clk),.wout(w76_92));
	PE pe76_93(.x(x93),.w(w76_92),.acc(r76_92),.res(r76_93),.clk(clk),.wout(w76_93));
	PE pe76_94(.x(x94),.w(w76_93),.acc(r76_93),.res(r76_94),.clk(clk),.wout(w76_94));
	PE pe76_95(.x(x95),.w(w76_94),.acc(r76_94),.res(r76_95),.clk(clk),.wout(w76_95));
	PE pe76_96(.x(x96),.w(w76_95),.acc(r76_95),.res(r76_96),.clk(clk),.wout(w76_96));
	PE pe76_97(.x(x97),.w(w76_96),.acc(r76_96),.res(r76_97),.clk(clk),.wout(w76_97));
	PE pe76_98(.x(x98),.w(w76_97),.acc(r76_97),.res(r76_98),.clk(clk),.wout(w76_98));
	PE pe76_99(.x(x99),.w(w76_98),.acc(r76_98),.res(r76_99),.clk(clk),.wout(w76_99));
	PE pe76_100(.x(x100),.w(w76_99),.acc(r76_99),.res(r76_100),.clk(clk),.wout(w76_100));
	PE pe76_101(.x(x101),.w(w76_100),.acc(r76_100),.res(r76_101),.clk(clk),.wout(w76_101));
	PE pe76_102(.x(x102),.w(w76_101),.acc(r76_101),.res(r76_102),.clk(clk),.wout(w76_102));
	PE pe76_103(.x(x103),.w(w76_102),.acc(r76_102),.res(r76_103),.clk(clk),.wout(w76_103));
	PE pe76_104(.x(x104),.w(w76_103),.acc(r76_103),.res(r76_104),.clk(clk),.wout(w76_104));
	PE pe76_105(.x(x105),.w(w76_104),.acc(r76_104),.res(r76_105),.clk(clk),.wout(w76_105));
	PE pe76_106(.x(x106),.w(w76_105),.acc(r76_105),.res(r76_106),.clk(clk),.wout(w76_106));
	PE pe76_107(.x(x107),.w(w76_106),.acc(r76_106),.res(r76_107),.clk(clk),.wout(w76_107));
	PE pe76_108(.x(x108),.w(w76_107),.acc(r76_107),.res(r76_108),.clk(clk),.wout(w76_108));
	PE pe76_109(.x(x109),.w(w76_108),.acc(r76_108),.res(r76_109),.clk(clk),.wout(w76_109));
	PE pe76_110(.x(x110),.w(w76_109),.acc(r76_109),.res(r76_110),.clk(clk),.wout(w76_110));
	PE pe76_111(.x(x111),.w(w76_110),.acc(r76_110),.res(r76_111),.clk(clk),.wout(w76_111));
	PE pe76_112(.x(x112),.w(w76_111),.acc(r76_111),.res(r76_112),.clk(clk),.wout(w76_112));
	PE pe76_113(.x(x113),.w(w76_112),.acc(r76_112),.res(r76_113),.clk(clk),.wout(w76_113));
	PE pe76_114(.x(x114),.w(w76_113),.acc(r76_113),.res(r76_114),.clk(clk),.wout(w76_114));
	PE pe76_115(.x(x115),.w(w76_114),.acc(r76_114),.res(r76_115),.clk(clk),.wout(w76_115));
	PE pe76_116(.x(x116),.w(w76_115),.acc(r76_115),.res(r76_116),.clk(clk),.wout(w76_116));
	PE pe76_117(.x(x117),.w(w76_116),.acc(r76_116),.res(r76_117),.clk(clk),.wout(w76_117));
	PE pe76_118(.x(x118),.w(w76_117),.acc(r76_117),.res(r76_118),.clk(clk),.wout(w76_118));
	PE pe76_119(.x(x119),.w(w76_118),.acc(r76_118),.res(r76_119),.clk(clk),.wout(w76_119));
	PE pe76_120(.x(x120),.w(w76_119),.acc(r76_119),.res(r76_120),.clk(clk),.wout(w76_120));
	PE pe76_121(.x(x121),.w(w76_120),.acc(r76_120),.res(r76_121),.clk(clk),.wout(w76_121));
	PE pe76_122(.x(x122),.w(w76_121),.acc(r76_121),.res(r76_122),.clk(clk),.wout(w76_122));
	PE pe76_123(.x(x123),.w(w76_122),.acc(r76_122),.res(r76_123),.clk(clk),.wout(w76_123));
	PE pe76_124(.x(x124),.w(w76_123),.acc(r76_123),.res(r76_124),.clk(clk),.wout(w76_124));
	PE pe76_125(.x(x125),.w(w76_124),.acc(r76_124),.res(r76_125),.clk(clk),.wout(w76_125));
	PE pe76_126(.x(x126),.w(w76_125),.acc(r76_125),.res(r76_126),.clk(clk),.wout(w76_126));
	PE pe76_127(.x(x127),.w(w76_126),.acc(r76_126),.res(result76),.clk(clk),.wout(weight76));

	PE pe77_0(.x(x0),.w(w77),.acc(32'h0),.res(r77_0),.clk(clk),.wout(w77_0));
	PE pe77_1(.x(x1),.w(w77_0),.acc(r77_0),.res(r77_1),.clk(clk),.wout(w77_1));
	PE pe77_2(.x(x2),.w(w77_1),.acc(r77_1),.res(r77_2),.clk(clk),.wout(w77_2));
	PE pe77_3(.x(x3),.w(w77_2),.acc(r77_2),.res(r77_3),.clk(clk),.wout(w77_3));
	PE pe77_4(.x(x4),.w(w77_3),.acc(r77_3),.res(r77_4),.clk(clk),.wout(w77_4));
	PE pe77_5(.x(x5),.w(w77_4),.acc(r77_4),.res(r77_5),.clk(clk),.wout(w77_5));
	PE pe77_6(.x(x6),.w(w77_5),.acc(r77_5),.res(r77_6),.clk(clk),.wout(w77_6));
	PE pe77_7(.x(x7),.w(w77_6),.acc(r77_6),.res(r77_7),.clk(clk),.wout(w77_7));
	PE pe77_8(.x(x8),.w(w77_7),.acc(r77_7),.res(r77_8),.clk(clk),.wout(w77_8));
	PE pe77_9(.x(x9),.w(w77_8),.acc(r77_8),.res(r77_9),.clk(clk),.wout(w77_9));
	PE pe77_10(.x(x10),.w(w77_9),.acc(r77_9),.res(r77_10),.clk(clk),.wout(w77_10));
	PE pe77_11(.x(x11),.w(w77_10),.acc(r77_10),.res(r77_11),.clk(clk),.wout(w77_11));
	PE pe77_12(.x(x12),.w(w77_11),.acc(r77_11),.res(r77_12),.clk(clk),.wout(w77_12));
	PE pe77_13(.x(x13),.w(w77_12),.acc(r77_12),.res(r77_13),.clk(clk),.wout(w77_13));
	PE pe77_14(.x(x14),.w(w77_13),.acc(r77_13),.res(r77_14),.clk(clk),.wout(w77_14));
	PE pe77_15(.x(x15),.w(w77_14),.acc(r77_14),.res(r77_15),.clk(clk),.wout(w77_15));
	PE pe77_16(.x(x16),.w(w77_15),.acc(r77_15),.res(r77_16),.clk(clk),.wout(w77_16));
	PE pe77_17(.x(x17),.w(w77_16),.acc(r77_16),.res(r77_17),.clk(clk),.wout(w77_17));
	PE pe77_18(.x(x18),.w(w77_17),.acc(r77_17),.res(r77_18),.clk(clk),.wout(w77_18));
	PE pe77_19(.x(x19),.w(w77_18),.acc(r77_18),.res(r77_19),.clk(clk),.wout(w77_19));
	PE pe77_20(.x(x20),.w(w77_19),.acc(r77_19),.res(r77_20),.clk(clk),.wout(w77_20));
	PE pe77_21(.x(x21),.w(w77_20),.acc(r77_20),.res(r77_21),.clk(clk),.wout(w77_21));
	PE pe77_22(.x(x22),.w(w77_21),.acc(r77_21),.res(r77_22),.clk(clk),.wout(w77_22));
	PE pe77_23(.x(x23),.w(w77_22),.acc(r77_22),.res(r77_23),.clk(clk),.wout(w77_23));
	PE pe77_24(.x(x24),.w(w77_23),.acc(r77_23),.res(r77_24),.clk(clk),.wout(w77_24));
	PE pe77_25(.x(x25),.w(w77_24),.acc(r77_24),.res(r77_25),.clk(clk),.wout(w77_25));
	PE pe77_26(.x(x26),.w(w77_25),.acc(r77_25),.res(r77_26),.clk(clk),.wout(w77_26));
	PE pe77_27(.x(x27),.w(w77_26),.acc(r77_26),.res(r77_27),.clk(clk),.wout(w77_27));
	PE pe77_28(.x(x28),.w(w77_27),.acc(r77_27),.res(r77_28),.clk(clk),.wout(w77_28));
	PE pe77_29(.x(x29),.w(w77_28),.acc(r77_28),.res(r77_29),.clk(clk),.wout(w77_29));
	PE pe77_30(.x(x30),.w(w77_29),.acc(r77_29),.res(r77_30),.clk(clk),.wout(w77_30));
	PE pe77_31(.x(x31),.w(w77_30),.acc(r77_30),.res(r77_31),.clk(clk),.wout(w77_31));
	PE pe77_32(.x(x32),.w(w77_31),.acc(r77_31),.res(r77_32),.clk(clk),.wout(w77_32));
	PE pe77_33(.x(x33),.w(w77_32),.acc(r77_32),.res(r77_33),.clk(clk),.wout(w77_33));
	PE pe77_34(.x(x34),.w(w77_33),.acc(r77_33),.res(r77_34),.clk(clk),.wout(w77_34));
	PE pe77_35(.x(x35),.w(w77_34),.acc(r77_34),.res(r77_35),.clk(clk),.wout(w77_35));
	PE pe77_36(.x(x36),.w(w77_35),.acc(r77_35),.res(r77_36),.clk(clk),.wout(w77_36));
	PE pe77_37(.x(x37),.w(w77_36),.acc(r77_36),.res(r77_37),.clk(clk),.wout(w77_37));
	PE pe77_38(.x(x38),.w(w77_37),.acc(r77_37),.res(r77_38),.clk(clk),.wout(w77_38));
	PE pe77_39(.x(x39),.w(w77_38),.acc(r77_38),.res(r77_39),.clk(clk),.wout(w77_39));
	PE pe77_40(.x(x40),.w(w77_39),.acc(r77_39),.res(r77_40),.clk(clk),.wout(w77_40));
	PE pe77_41(.x(x41),.w(w77_40),.acc(r77_40),.res(r77_41),.clk(clk),.wout(w77_41));
	PE pe77_42(.x(x42),.w(w77_41),.acc(r77_41),.res(r77_42),.clk(clk),.wout(w77_42));
	PE pe77_43(.x(x43),.w(w77_42),.acc(r77_42),.res(r77_43),.clk(clk),.wout(w77_43));
	PE pe77_44(.x(x44),.w(w77_43),.acc(r77_43),.res(r77_44),.clk(clk),.wout(w77_44));
	PE pe77_45(.x(x45),.w(w77_44),.acc(r77_44),.res(r77_45),.clk(clk),.wout(w77_45));
	PE pe77_46(.x(x46),.w(w77_45),.acc(r77_45),.res(r77_46),.clk(clk),.wout(w77_46));
	PE pe77_47(.x(x47),.w(w77_46),.acc(r77_46),.res(r77_47),.clk(clk),.wout(w77_47));
	PE pe77_48(.x(x48),.w(w77_47),.acc(r77_47),.res(r77_48),.clk(clk),.wout(w77_48));
	PE pe77_49(.x(x49),.w(w77_48),.acc(r77_48),.res(r77_49),.clk(clk),.wout(w77_49));
	PE pe77_50(.x(x50),.w(w77_49),.acc(r77_49),.res(r77_50),.clk(clk),.wout(w77_50));
	PE pe77_51(.x(x51),.w(w77_50),.acc(r77_50),.res(r77_51),.clk(clk),.wout(w77_51));
	PE pe77_52(.x(x52),.w(w77_51),.acc(r77_51),.res(r77_52),.clk(clk),.wout(w77_52));
	PE pe77_53(.x(x53),.w(w77_52),.acc(r77_52),.res(r77_53),.clk(clk),.wout(w77_53));
	PE pe77_54(.x(x54),.w(w77_53),.acc(r77_53),.res(r77_54),.clk(clk),.wout(w77_54));
	PE pe77_55(.x(x55),.w(w77_54),.acc(r77_54),.res(r77_55),.clk(clk),.wout(w77_55));
	PE pe77_56(.x(x56),.w(w77_55),.acc(r77_55),.res(r77_56),.clk(clk),.wout(w77_56));
	PE pe77_57(.x(x57),.w(w77_56),.acc(r77_56),.res(r77_57),.clk(clk),.wout(w77_57));
	PE pe77_58(.x(x58),.w(w77_57),.acc(r77_57),.res(r77_58),.clk(clk),.wout(w77_58));
	PE pe77_59(.x(x59),.w(w77_58),.acc(r77_58),.res(r77_59),.clk(clk),.wout(w77_59));
	PE pe77_60(.x(x60),.w(w77_59),.acc(r77_59),.res(r77_60),.clk(clk),.wout(w77_60));
	PE pe77_61(.x(x61),.w(w77_60),.acc(r77_60),.res(r77_61),.clk(clk),.wout(w77_61));
	PE pe77_62(.x(x62),.w(w77_61),.acc(r77_61),.res(r77_62),.clk(clk),.wout(w77_62));
	PE pe77_63(.x(x63),.w(w77_62),.acc(r77_62),.res(r77_63),.clk(clk),.wout(w77_63));
	PE pe77_64(.x(x64),.w(w77_63),.acc(r77_63),.res(r77_64),.clk(clk),.wout(w77_64));
	PE pe77_65(.x(x65),.w(w77_64),.acc(r77_64),.res(r77_65),.clk(clk),.wout(w77_65));
	PE pe77_66(.x(x66),.w(w77_65),.acc(r77_65),.res(r77_66),.clk(clk),.wout(w77_66));
	PE pe77_67(.x(x67),.w(w77_66),.acc(r77_66),.res(r77_67),.clk(clk),.wout(w77_67));
	PE pe77_68(.x(x68),.w(w77_67),.acc(r77_67),.res(r77_68),.clk(clk),.wout(w77_68));
	PE pe77_69(.x(x69),.w(w77_68),.acc(r77_68),.res(r77_69),.clk(clk),.wout(w77_69));
	PE pe77_70(.x(x70),.w(w77_69),.acc(r77_69),.res(r77_70),.clk(clk),.wout(w77_70));
	PE pe77_71(.x(x71),.w(w77_70),.acc(r77_70),.res(r77_71),.clk(clk),.wout(w77_71));
	PE pe77_72(.x(x72),.w(w77_71),.acc(r77_71),.res(r77_72),.clk(clk),.wout(w77_72));
	PE pe77_73(.x(x73),.w(w77_72),.acc(r77_72),.res(r77_73),.clk(clk),.wout(w77_73));
	PE pe77_74(.x(x74),.w(w77_73),.acc(r77_73),.res(r77_74),.clk(clk),.wout(w77_74));
	PE pe77_75(.x(x75),.w(w77_74),.acc(r77_74),.res(r77_75),.clk(clk),.wout(w77_75));
	PE pe77_76(.x(x76),.w(w77_75),.acc(r77_75),.res(r77_76),.clk(clk),.wout(w77_76));
	PE pe77_77(.x(x77),.w(w77_76),.acc(r77_76),.res(r77_77),.clk(clk),.wout(w77_77));
	PE pe77_78(.x(x78),.w(w77_77),.acc(r77_77),.res(r77_78),.clk(clk),.wout(w77_78));
	PE pe77_79(.x(x79),.w(w77_78),.acc(r77_78),.res(r77_79),.clk(clk),.wout(w77_79));
	PE pe77_80(.x(x80),.w(w77_79),.acc(r77_79),.res(r77_80),.clk(clk),.wout(w77_80));
	PE pe77_81(.x(x81),.w(w77_80),.acc(r77_80),.res(r77_81),.clk(clk),.wout(w77_81));
	PE pe77_82(.x(x82),.w(w77_81),.acc(r77_81),.res(r77_82),.clk(clk),.wout(w77_82));
	PE pe77_83(.x(x83),.w(w77_82),.acc(r77_82),.res(r77_83),.clk(clk),.wout(w77_83));
	PE pe77_84(.x(x84),.w(w77_83),.acc(r77_83),.res(r77_84),.clk(clk),.wout(w77_84));
	PE pe77_85(.x(x85),.w(w77_84),.acc(r77_84),.res(r77_85),.clk(clk),.wout(w77_85));
	PE pe77_86(.x(x86),.w(w77_85),.acc(r77_85),.res(r77_86),.clk(clk),.wout(w77_86));
	PE pe77_87(.x(x87),.w(w77_86),.acc(r77_86),.res(r77_87),.clk(clk),.wout(w77_87));
	PE pe77_88(.x(x88),.w(w77_87),.acc(r77_87),.res(r77_88),.clk(clk),.wout(w77_88));
	PE pe77_89(.x(x89),.w(w77_88),.acc(r77_88),.res(r77_89),.clk(clk),.wout(w77_89));
	PE pe77_90(.x(x90),.w(w77_89),.acc(r77_89),.res(r77_90),.clk(clk),.wout(w77_90));
	PE pe77_91(.x(x91),.w(w77_90),.acc(r77_90),.res(r77_91),.clk(clk),.wout(w77_91));
	PE pe77_92(.x(x92),.w(w77_91),.acc(r77_91),.res(r77_92),.clk(clk),.wout(w77_92));
	PE pe77_93(.x(x93),.w(w77_92),.acc(r77_92),.res(r77_93),.clk(clk),.wout(w77_93));
	PE pe77_94(.x(x94),.w(w77_93),.acc(r77_93),.res(r77_94),.clk(clk),.wout(w77_94));
	PE pe77_95(.x(x95),.w(w77_94),.acc(r77_94),.res(r77_95),.clk(clk),.wout(w77_95));
	PE pe77_96(.x(x96),.w(w77_95),.acc(r77_95),.res(r77_96),.clk(clk),.wout(w77_96));
	PE pe77_97(.x(x97),.w(w77_96),.acc(r77_96),.res(r77_97),.clk(clk),.wout(w77_97));
	PE pe77_98(.x(x98),.w(w77_97),.acc(r77_97),.res(r77_98),.clk(clk),.wout(w77_98));
	PE pe77_99(.x(x99),.w(w77_98),.acc(r77_98),.res(r77_99),.clk(clk),.wout(w77_99));
	PE pe77_100(.x(x100),.w(w77_99),.acc(r77_99),.res(r77_100),.clk(clk),.wout(w77_100));
	PE pe77_101(.x(x101),.w(w77_100),.acc(r77_100),.res(r77_101),.clk(clk),.wout(w77_101));
	PE pe77_102(.x(x102),.w(w77_101),.acc(r77_101),.res(r77_102),.clk(clk),.wout(w77_102));
	PE pe77_103(.x(x103),.w(w77_102),.acc(r77_102),.res(r77_103),.clk(clk),.wout(w77_103));
	PE pe77_104(.x(x104),.w(w77_103),.acc(r77_103),.res(r77_104),.clk(clk),.wout(w77_104));
	PE pe77_105(.x(x105),.w(w77_104),.acc(r77_104),.res(r77_105),.clk(clk),.wout(w77_105));
	PE pe77_106(.x(x106),.w(w77_105),.acc(r77_105),.res(r77_106),.clk(clk),.wout(w77_106));
	PE pe77_107(.x(x107),.w(w77_106),.acc(r77_106),.res(r77_107),.clk(clk),.wout(w77_107));
	PE pe77_108(.x(x108),.w(w77_107),.acc(r77_107),.res(r77_108),.clk(clk),.wout(w77_108));
	PE pe77_109(.x(x109),.w(w77_108),.acc(r77_108),.res(r77_109),.clk(clk),.wout(w77_109));
	PE pe77_110(.x(x110),.w(w77_109),.acc(r77_109),.res(r77_110),.clk(clk),.wout(w77_110));
	PE pe77_111(.x(x111),.w(w77_110),.acc(r77_110),.res(r77_111),.clk(clk),.wout(w77_111));
	PE pe77_112(.x(x112),.w(w77_111),.acc(r77_111),.res(r77_112),.clk(clk),.wout(w77_112));
	PE pe77_113(.x(x113),.w(w77_112),.acc(r77_112),.res(r77_113),.clk(clk),.wout(w77_113));
	PE pe77_114(.x(x114),.w(w77_113),.acc(r77_113),.res(r77_114),.clk(clk),.wout(w77_114));
	PE pe77_115(.x(x115),.w(w77_114),.acc(r77_114),.res(r77_115),.clk(clk),.wout(w77_115));
	PE pe77_116(.x(x116),.w(w77_115),.acc(r77_115),.res(r77_116),.clk(clk),.wout(w77_116));
	PE pe77_117(.x(x117),.w(w77_116),.acc(r77_116),.res(r77_117),.clk(clk),.wout(w77_117));
	PE pe77_118(.x(x118),.w(w77_117),.acc(r77_117),.res(r77_118),.clk(clk),.wout(w77_118));
	PE pe77_119(.x(x119),.w(w77_118),.acc(r77_118),.res(r77_119),.clk(clk),.wout(w77_119));
	PE pe77_120(.x(x120),.w(w77_119),.acc(r77_119),.res(r77_120),.clk(clk),.wout(w77_120));
	PE pe77_121(.x(x121),.w(w77_120),.acc(r77_120),.res(r77_121),.clk(clk),.wout(w77_121));
	PE pe77_122(.x(x122),.w(w77_121),.acc(r77_121),.res(r77_122),.clk(clk),.wout(w77_122));
	PE pe77_123(.x(x123),.w(w77_122),.acc(r77_122),.res(r77_123),.clk(clk),.wout(w77_123));
	PE pe77_124(.x(x124),.w(w77_123),.acc(r77_123),.res(r77_124),.clk(clk),.wout(w77_124));
	PE pe77_125(.x(x125),.w(w77_124),.acc(r77_124),.res(r77_125),.clk(clk),.wout(w77_125));
	PE pe77_126(.x(x126),.w(w77_125),.acc(r77_125),.res(r77_126),.clk(clk),.wout(w77_126));
	PE pe77_127(.x(x127),.w(w77_126),.acc(r77_126),.res(result77),.clk(clk),.wout(weight77));

	PE pe78_0(.x(x0),.w(w78),.acc(32'h0),.res(r78_0),.clk(clk),.wout(w78_0));
	PE pe78_1(.x(x1),.w(w78_0),.acc(r78_0),.res(r78_1),.clk(clk),.wout(w78_1));
	PE pe78_2(.x(x2),.w(w78_1),.acc(r78_1),.res(r78_2),.clk(clk),.wout(w78_2));
	PE pe78_3(.x(x3),.w(w78_2),.acc(r78_2),.res(r78_3),.clk(clk),.wout(w78_3));
	PE pe78_4(.x(x4),.w(w78_3),.acc(r78_3),.res(r78_4),.clk(clk),.wout(w78_4));
	PE pe78_5(.x(x5),.w(w78_4),.acc(r78_4),.res(r78_5),.clk(clk),.wout(w78_5));
	PE pe78_6(.x(x6),.w(w78_5),.acc(r78_5),.res(r78_6),.clk(clk),.wout(w78_6));
	PE pe78_7(.x(x7),.w(w78_6),.acc(r78_6),.res(r78_7),.clk(clk),.wout(w78_7));
	PE pe78_8(.x(x8),.w(w78_7),.acc(r78_7),.res(r78_8),.clk(clk),.wout(w78_8));
	PE pe78_9(.x(x9),.w(w78_8),.acc(r78_8),.res(r78_9),.clk(clk),.wout(w78_9));
	PE pe78_10(.x(x10),.w(w78_9),.acc(r78_9),.res(r78_10),.clk(clk),.wout(w78_10));
	PE pe78_11(.x(x11),.w(w78_10),.acc(r78_10),.res(r78_11),.clk(clk),.wout(w78_11));
	PE pe78_12(.x(x12),.w(w78_11),.acc(r78_11),.res(r78_12),.clk(clk),.wout(w78_12));
	PE pe78_13(.x(x13),.w(w78_12),.acc(r78_12),.res(r78_13),.clk(clk),.wout(w78_13));
	PE pe78_14(.x(x14),.w(w78_13),.acc(r78_13),.res(r78_14),.clk(clk),.wout(w78_14));
	PE pe78_15(.x(x15),.w(w78_14),.acc(r78_14),.res(r78_15),.clk(clk),.wout(w78_15));
	PE pe78_16(.x(x16),.w(w78_15),.acc(r78_15),.res(r78_16),.clk(clk),.wout(w78_16));
	PE pe78_17(.x(x17),.w(w78_16),.acc(r78_16),.res(r78_17),.clk(clk),.wout(w78_17));
	PE pe78_18(.x(x18),.w(w78_17),.acc(r78_17),.res(r78_18),.clk(clk),.wout(w78_18));
	PE pe78_19(.x(x19),.w(w78_18),.acc(r78_18),.res(r78_19),.clk(clk),.wout(w78_19));
	PE pe78_20(.x(x20),.w(w78_19),.acc(r78_19),.res(r78_20),.clk(clk),.wout(w78_20));
	PE pe78_21(.x(x21),.w(w78_20),.acc(r78_20),.res(r78_21),.clk(clk),.wout(w78_21));
	PE pe78_22(.x(x22),.w(w78_21),.acc(r78_21),.res(r78_22),.clk(clk),.wout(w78_22));
	PE pe78_23(.x(x23),.w(w78_22),.acc(r78_22),.res(r78_23),.clk(clk),.wout(w78_23));
	PE pe78_24(.x(x24),.w(w78_23),.acc(r78_23),.res(r78_24),.clk(clk),.wout(w78_24));
	PE pe78_25(.x(x25),.w(w78_24),.acc(r78_24),.res(r78_25),.clk(clk),.wout(w78_25));
	PE pe78_26(.x(x26),.w(w78_25),.acc(r78_25),.res(r78_26),.clk(clk),.wout(w78_26));
	PE pe78_27(.x(x27),.w(w78_26),.acc(r78_26),.res(r78_27),.clk(clk),.wout(w78_27));
	PE pe78_28(.x(x28),.w(w78_27),.acc(r78_27),.res(r78_28),.clk(clk),.wout(w78_28));
	PE pe78_29(.x(x29),.w(w78_28),.acc(r78_28),.res(r78_29),.clk(clk),.wout(w78_29));
	PE pe78_30(.x(x30),.w(w78_29),.acc(r78_29),.res(r78_30),.clk(clk),.wout(w78_30));
	PE pe78_31(.x(x31),.w(w78_30),.acc(r78_30),.res(r78_31),.clk(clk),.wout(w78_31));
	PE pe78_32(.x(x32),.w(w78_31),.acc(r78_31),.res(r78_32),.clk(clk),.wout(w78_32));
	PE pe78_33(.x(x33),.w(w78_32),.acc(r78_32),.res(r78_33),.clk(clk),.wout(w78_33));
	PE pe78_34(.x(x34),.w(w78_33),.acc(r78_33),.res(r78_34),.clk(clk),.wout(w78_34));
	PE pe78_35(.x(x35),.w(w78_34),.acc(r78_34),.res(r78_35),.clk(clk),.wout(w78_35));
	PE pe78_36(.x(x36),.w(w78_35),.acc(r78_35),.res(r78_36),.clk(clk),.wout(w78_36));
	PE pe78_37(.x(x37),.w(w78_36),.acc(r78_36),.res(r78_37),.clk(clk),.wout(w78_37));
	PE pe78_38(.x(x38),.w(w78_37),.acc(r78_37),.res(r78_38),.clk(clk),.wout(w78_38));
	PE pe78_39(.x(x39),.w(w78_38),.acc(r78_38),.res(r78_39),.clk(clk),.wout(w78_39));
	PE pe78_40(.x(x40),.w(w78_39),.acc(r78_39),.res(r78_40),.clk(clk),.wout(w78_40));
	PE pe78_41(.x(x41),.w(w78_40),.acc(r78_40),.res(r78_41),.clk(clk),.wout(w78_41));
	PE pe78_42(.x(x42),.w(w78_41),.acc(r78_41),.res(r78_42),.clk(clk),.wout(w78_42));
	PE pe78_43(.x(x43),.w(w78_42),.acc(r78_42),.res(r78_43),.clk(clk),.wout(w78_43));
	PE pe78_44(.x(x44),.w(w78_43),.acc(r78_43),.res(r78_44),.clk(clk),.wout(w78_44));
	PE pe78_45(.x(x45),.w(w78_44),.acc(r78_44),.res(r78_45),.clk(clk),.wout(w78_45));
	PE pe78_46(.x(x46),.w(w78_45),.acc(r78_45),.res(r78_46),.clk(clk),.wout(w78_46));
	PE pe78_47(.x(x47),.w(w78_46),.acc(r78_46),.res(r78_47),.clk(clk),.wout(w78_47));
	PE pe78_48(.x(x48),.w(w78_47),.acc(r78_47),.res(r78_48),.clk(clk),.wout(w78_48));
	PE pe78_49(.x(x49),.w(w78_48),.acc(r78_48),.res(r78_49),.clk(clk),.wout(w78_49));
	PE pe78_50(.x(x50),.w(w78_49),.acc(r78_49),.res(r78_50),.clk(clk),.wout(w78_50));
	PE pe78_51(.x(x51),.w(w78_50),.acc(r78_50),.res(r78_51),.clk(clk),.wout(w78_51));
	PE pe78_52(.x(x52),.w(w78_51),.acc(r78_51),.res(r78_52),.clk(clk),.wout(w78_52));
	PE pe78_53(.x(x53),.w(w78_52),.acc(r78_52),.res(r78_53),.clk(clk),.wout(w78_53));
	PE pe78_54(.x(x54),.w(w78_53),.acc(r78_53),.res(r78_54),.clk(clk),.wout(w78_54));
	PE pe78_55(.x(x55),.w(w78_54),.acc(r78_54),.res(r78_55),.clk(clk),.wout(w78_55));
	PE pe78_56(.x(x56),.w(w78_55),.acc(r78_55),.res(r78_56),.clk(clk),.wout(w78_56));
	PE pe78_57(.x(x57),.w(w78_56),.acc(r78_56),.res(r78_57),.clk(clk),.wout(w78_57));
	PE pe78_58(.x(x58),.w(w78_57),.acc(r78_57),.res(r78_58),.clk(clk),.wout(w78_58));
	PE pe78_59(.x(x59),.w(w78_58),.acc(r78_58),.res(r78_59),.clk(clk),.wout(w78_59));
	PE pe78_60(.x(x60),.w(w78_59),.acc(r78_59),.res(r78_60),.clk(clk),.wout(w78_60));
	PE pe78_61(.x(x61),.w(w78_60),.acc(r78_60),.res(r78_61),.clk(clk),.wout(w78_61));
	PE pe78_62(.x(x62),.w(w78_61),.acc(r78_61),.res(r78_62),.clk(clk),.wout(w78_62));
	PE pe78_63(.x(x63),.w(w78_62),.acc(r78_62),.res(r78_63),.clk(clk),.wout(w78_63));
	PE pe78_64(.x(x64),.w(w78_63),.acc(r78_63),.res(r78_64),.clk(clk),.wout(w78_64));
	PE pe78_65(.x(x65),.w(w78_64),.acc(r78_64),.res(r78_65),.clk(clk),.wout(w78_65));
	PE pe78_66(.x(x66),.w(w78_65),.acc(r78_65),.res(r78_66),.clk(clk),.wout(w78_66));
	PE pe78_67(.x(x67),.w(w78_66),.acc(r78_66),.res(r78_67),.clk(clk),.wout(w78_67));
	PE pe78_68(.x(x68),.w(w78_67),.acc(r78_67),.res(r78_68),.clk(clk),.wout(w78_68));
	PE pe78_69(.x(x69),.w(w78_68),.acc(r78_68),.res(r78_69),.clk(clk),.wout(w78_69));
	PE pe78_70(.x(x70),.w(w78_69),.acc(r78_69),.res(r78_70),.clk(clk),.wout(w78_70));
	PE pe78_71(.x(x71),.w(w78_70),.acc(r78_70),.res(r78_71),.clk(clk),.wout(w78_71));
	PE pe78_72(.x(x72),.w(w78_71),.acc(r78_71),.res(r78_72),.clk(clk),.wout(w78_72));
	PE pe78_73(.x(x73),.w(w78_72),.acc(r78_72),.res(r78_73),.clk(clk),.wout(w78_73));
	PE pe78_74(.x(x74),.w(w78_73),.acc(r78_73),.res(r78_74),.clk(clk),.wout(w78_74));
	PE pe78_75(.x(x75),.w(w78_74),.acc(r78_74),.res(r78_75),.clk(clk),.wout(w78_75));
	PE pe78_76(.x(x76),.w(w78_75),.acc(r78_75),.res(r78_76),.clk(clk),.wout(w78_76));
	PE pe78_77(.x(x77),.w(w78_76),.acc(r78_76),.res(r78_77),.clk(clk),.wout(w78_77));
	PE pe78_78(.x(x78),.w(w78_77),.acc(r78_77),.res(r78_78),.clk(clk),.wout(w78_78));
	PE pe78_79(.x(x79),.w(w78_78),.acc(r78_78),.res(r78_79),.clk(clk),.wout(w78_79));
	PE pe78_80(.x(x80),.w(w78_79),.acc(r78_79),.res(r78_80),.clk(clk),.wout(w78_80));
	PE pe78_81(.x(x81),.w(w78_80),.acc(r78_80),.res(r78_81),.clk(clk),.wout(w78_81));
	PE pe78_82(.x(x82),.w(w78_81),.acc(r78_81),.res(r78_82),.clk(clk),.wout(w78_82));
	PE pe78_83(.x(x83),.w(w78_82),.acc(r78_82),.res(r78_83),.clk(clk),.wout(w78_83));
	PE pe78_84(.x(x84),.w(w78_83),.acc(r78_83),.res(r78_84),.clk(clk),.wout(w78_84));
	PE pe78_85(.x(x85),.w(w78_84),.acc(r78_84),.res(r78_85),.clk(clk),.wout(w78_85));
	PE pe78_86(.x(x86),.w(w78_85),.acc(r78_85),.res(r78_86),.clk(clk),.wout(w78_86));
	PE pe78_87(.x(x87),.w(w78_86),.acc(r78_86),.res(r78_87),.clk(clk),.wout(w78_87));
	PE pe78_88(.x(x88),.w(w78_87),.acc(r78_87),.res(r78_88),.clk(clk),.wout(w78_88));
	PE pe78_89(.x(x89),.w(w78_88),.acc(r78_88),.res(r78_89),.clk(clk),.wout(w78_89));
	PE pe78_90(.x(x90),.w(w78_89),.acc(r78_89),.res(r78_90),.clk(clk),.wout(w78_90));
	PE pe78_91(.x(x91),.w(w78_90),.acc(r78_90),.res(r78_91),.clk(clk),.wout(w78_91));
	PE pe78_92(.x(x92),.w(w78_91),.acc(r78_91),.res(r78_92),.clk(clk),.wout(w78_92));
	PE pe78_93(.x(x93),.w(w78_92),.acc(r78_92),.res(r78_93),.clk(clk),.wout(w78_93));
	PE pe78_94(.x(x94),.w(w78_93),.acc(r78_93),.res(r78_94),.clk(clk),.wout(w78_94));
	PE pe78_95(.x(x95),.w(w78_94),.acc(r78_94),.res(r78_95),.clk(clk),.wout(w78_95));
	PE pe78_96(.x(x96),.w(w78_95),.acc(r78_95),.res(r78_96),.clk(clk),.wout(w78_96));
	PE pe78_97(.x(x97),.w(w78_96),.acc(r78_96),.res(r78_97),.clk(clk),.wout(w78_97));
	PE pe78_98(.x(x98),.w(w78_97),.acc(r78_97),.res(r78_98),.clk(clk),.wout(w78_98));
	PE pe78_99(.x(x99),.w(w78_98),.acc(r78_98),.res(r78_99),.clk(clk),.wout(w78_99));
	PE pe78_100(.x(x100),.w(w78_99),.acc(r78_99),.res(r78_100),.clk(clk),.wout(w78_100));
	PE pe78_101(.x(x101),.w(w78_100),.acc(r78_100),.res(r78_101),.clk(clk),.wout(w78_101));
	PE pe78_102(.x(x102),.w(w78_101),.acc(r78_101),.res(r78_102),.clk(clk),.wout(w78_102));
	PE pe78_103(.x(x103),.w(w78_102),.acc(r78_102),.res(r78_103),.clk(clk),.wout(w78_103));
	PE pe78_104(.x(x104),.w(w78_103),.acc(r78_103),.res(r78_104),.clk(clk),.wout(w78_104));
	PE pe78_105(.x(x105),.w(w78_104),.acc(r78_104),.res(r78_105),.clk(clk),.wout(w78_105));
	PE pe78_106(.x(x106),.w(w78_105),.acc(r78_105),.res(r78_106),.clk(clk),.wout(w78_106));
	PE pe78_107(.x(x107),.w(w78_106),.acc(r78_106),.res(r78_107),.clk(clk),.wout(w78_107));
	PE pe78_108(.x(x108),.w(w78_107),.acc(r78_107),.res(r78_108),.clk(clk),.wout(w78_108));
	PE pe78_109(.x(x109),.w(w78_108),.acc(r78_108),.res(r78_109),.clk(clk),.wout(w78_109));
	PE pe78_110(.x(x110),.w(w78_109),.acc(r78_109),.res(r78_110),.clk(clk),.wout(w78_110));
	PE pe78_111(.x(x111),.w(w78_110),.acc(r78_110),.res(r78_111),.clk(clk),.wout(w78_111));
	PE pe78_112(.x(x112),.w(w78_111),.acc(r78_111),.res(r78_112),.clk(clk),.wout(w78_112));
	PE pe78_113(.x(x113),.w(w78_112),.acc(r78_112),.res(r78_113),.clk(clk),.wout(w78_113));
	PE pe78_114(.x(x114),.w(w78_113),.acc(r78_113),.res(r78_114),.clk(clk),.wout(w78_114));
	PE pe78_115(.x(x115),.w(w78_114),.acc(r78_114),.res(r78_115),.clk(clk),.wout(w78_115));
	PE pe78_116(.x(x116),.w(w78_115),.acc(r78_115),.res(r78_116),.clk(clk),.wout(w78_116));
	PE pe78_117(.x(x117),.w(w78_116),.acc(r78_116),.res(r78_117),.clk(clk),.wout(w78_117));
	PE pe78_118(.x(x118),.w(w78_117),.acc(r78_117),.res(r78_118),.clk(clk),.wout(w78_118));
	PE pe78_119(.x(x119),.w(w78_118),.acc(r78_118),.res(r78_119),.clk(clk),.wout(w78_119));
	PE pe78_120(.x(x120),.w(w78_119),.acc(r78_119),.res(r78_120),.clk(clk),.wout(w78_120));
	PE pe78_121(.x(x121),.w(w78_120),.acc(r78_120),.res(r78_121),.clk(clk),.wout(w78_121));
	PE pe78_122(.x(x122),.w(w78_121),.acc(r78_121),.res(r78_122),.clk(clk),.wout(w78_122));
	PE pe78_123(.x(x123),.w(w78_122),.acc(r78_122),.res(r78_123),.clk(clk),.wout(w78_123));
	PE pe78_124(.x(x124),.w(w78_123),.acc(r78_123),.res(r78_124),.clk(clk),.wout(w78_124));
	PE pe78_125(.x(x125),.w(w78_124),.acc(r78_124),.res(r78_125),.clk(clk),.wout(w78_125));
	PE pe78_126(.x(x126),.w(w78_125),.acc(r78_125),.res(r78_126),.clk(clk),.wout(w78_126));
	PE pe78_127(.x(x127),.w(w78_126),.acc(r78_126),.res(result78),.clk(clk),.wout(weight78));

	PE pe79_0(.x(x0),.w(w79),.acc(32'h0),.res(r79_0),.clk(clk),.wout(w79_0));
	PE pe79_1(.x(x1),.w(w79_0),.acc(r79_0),.res(r79_1),.clk(clk),.wout(w79_1));
	PE pe79_2(.x(x2),.w(w79_1),.acc(r79_1),.res(r79_2),.clk(clk),.wout(w79_2));
	PE pe79_3(.x(x3),.w(w79_2),.acc(r79_2),.res(r79_3),.clk(clk),.wout(w79_3));
	PE pe79_4(.x(x4),.w(w79_3),.acc(r79_3),.res(r79_4),.clk(clk),.wout(w79_4));
	PE pe79_5(.x(x5),.w(w79_4),.acc(r79_4),.res(r79_5),.clk(clk),.wout(w79_5));
	PE pe79_6(.x(x6),.w(w79_5),.acc(r79_5),.res(r79_6),.clk(clk),.wout(w79_6));
	PE pe79_7(.x(x7),.w(w79_6),.acc(r79_6),.res(r79_7),.clk(clk),.wout(w79_7));
	PE pe79_8(.x(x8),.w(w79_7),.acc(r79_7),.res(r79_8),.clk(clk),.wout(w79_8));
	PE pe79_9(.x(x9),.w(w79_8),.acc(r79_8),.res(r79_9),.clk(clk),.wout(w79_9));
	PE pe79_10(.x(x10),.w(w79_9),.acc(r79_9),.res(r79_10),.clk(clk),.wout(w79_10));
	PE pe79_11(.x(x11),.w(w79_10),.acc(r79_10),.res(r79_11),.clk(clk),.wout(w79_11));
	PE pe79_12(.x(x12),.w(w79_11),.acc(r79_11),.res(r79_12),.clk(clk),.wout(w79_12));
	PE pe79_13(.x(x13),.w(w79_12),.acc(r79_12),.res(r79_13),.clk(clk),.wout(w79_13));
	PE pe79_14(.x(x14),.w(w79_13),.acc(r79_13),.res(r79_14),.clk(clk),.wout(w79_14));
	PE pe79_15(.x(x15),.w(w79_14),.acc(r79_14),.res(r79_15),.clk(clk),.wout(w79_15));
	PE pe79_16(.x(x16),.w(w79_15),.acc(r79_15),.res(r79_16),.clk(clk),.wout(w79_16));
	PE pe79_17(.x(x17),.w(w79_16),.acc(r79_16),.res(r79_17),.clk(clk),.wout(w79_17));
	PE pe79_18(.x(x18),.w(w79_17),.acc(r79_17),.res(r79_18),.clk(clk),.wout(w79_18));
	PE pe79_19(.x(x19),.w(w79_18),.acc(r79_18),.res(r79_19),.clk(clk),.wout(w79_19));
	PE pe79_20(.x(x20),.w(w79_19),.acc(r79_19),.res(r79_20),.clk(clk),.wout(w79_20));
	PE pe79_21(.x(x21),.w(w79_20),.acc(r79_20),.res(r79_21),.clk(clk),.wout(w79_21));
	PE pe79_22(.x(x22),.w(w79_21),.acc(r79_21),.res(r79_22),.clk(clk),.wout(w79_22));
	PE pe79_23(.x(x23),.w(w79_22),.acc(r79_22),.res(r79_23),.clk(clk),.wout(w79_23));
	PE pe79_24(.x(x24),.w(w79_23),.acc(r79_23),.res(r79_24),.clk(clk),.wout(w79_24));
	PE pe79_25(.x(x25),.w(w79_24),.acc(r79_24),.res(r79_25),.clk(clk),.wout(w79_25));
	PE pe79_26(.x(x26),.w(w79_25),.acc(r79_25),.res(r79_26),.clk(clk),.wout(w79_26));
	PE pe79_27(.x(x27),.w(w79_26),.acc(r79_26),.res(r79_27),.clk(clk),.wout(w79_27));
	PE pe79_28(.x(x28),.w(w79_27),.acc(r79_27),.res(r79_28),.clk(clk),.wout(w79_28));
	PE pe79_29(.x(x29),.w(w79_28),.acc(r79_28),.res(r79_29),.clk(clk),.wout(w79_29));
	PE pe79_30(.x(x30),.w(w79_29),.acc(r79_29),.res(r79_30),.clk(clk),.wout(w79_30));
	PE pe79_31(.x(x31),.w(w79_30),.acc(r79_30),.res(r79_31),.clk(clk),.wout(w79_31));
	PE pe79_32(.x(x32),.w(w79_31),.acc(r79_31),.res(r79_32),.clk(clk),.wout(w79_32));
	PE pe79_33(.x(x33),.w(w79_32),.acc(r79_32),.res(r79_33),.clk(clk),.wout(w79_33));
	PE pe79_34(.x(x34),.w(w79_33),.acc(r79_33),.res(r79_34),.clk(clk),.wout(w79_34));
	PE pe79_35(.x(x35),.w(w79_34),.acc(r79_34),.res(r79_35),.clk(clk),.wout(w79_35));
	PE pe79_36(.x(x36),.w(w79_35),.acc(r79_35),.res(r79_36),.clk(clk),.wout(w79_36));
	PE pe79_37(.x(x37),.w(w79_36),.acc(r79_36),.res(r79_37),.clk(clk),.wout(w79_37));
	PE pe79_38(.x(x38),.w(w79_37),.acc(r79_37),.res(r79_38),.clk(clk),.wout(w79_38));
	PE pe79_39(.x(x39),.w(w79_38),.acc(r79_38),.res(r79_39),.clk(clk),.wout(w79_39));
	PE pe79_40(.x(x40),.w(w79_39),.acc(r79_39),.res(r79_40),.clk(clk),.wout(w79_40));
	PE pe79_41(.x(x41),.w(w79_40),.acc(r79_40),.res(r79_41),.clk(clk),.wout(w79_41));
	PE pe79_42(.x(x42),.w(w79_41),.acc(r79_41),.res(r79_42),.clk(clk),.wout(w79_42));
	PE pe79_43(.x(x43),.w(w79_42),.acc(r79_42),.res(r79_43),.clk(clk),.wout(w79_43));
	PE pe79_44(.x(x44),.w(w79_43),.acc(r79_43),.res(r79_44),.clk(clk),.wout(w79_44));
	PE pe79_45(.x(x45),.w(w79_44),.acc(r79_44),.res(r79_45),.clk(clk),.wout(w79_45));
	PE pe79_46(.x(x46),.w(w79_45),.acc(r79_45),.res(r79_46),.clk(clk),.wout(w79_46));
	PE pe79_47(.x(x47),.w(w79_46),.acc(r79_46),.res(r79_47),.clk(clk),.wout(w79_47));
	PE pe79_48(.x(x48),.w(w79_47),.acc(r79_47),.res(r79_48),.clk(clk),.wout(w79_48));
	PE pe79_49(.x(x49),.w(w79_48),.acc(r79_48),.res(r79_49),.clk(clk),.wout(w79_49));
	PE pe79_50(.x(x50),.w(w79_49),.acc(r79_49),.res(r79_50),.clk(clk),.wout(w79_50));
	PE pe79_51(.x(x51),.w(w79_50),.acc(r79_50),.res(r79_51),.clk(clk),.wout(w79_51));
	PE pe79_52(.x(x52),.w(w79_51),.acc(r79_51),.res(r79_52),.clk(clk),.wout(w79_52));
	PE pe79_53(.x(x53),.w(w79_52),.acc(r79_52),.res(r79_53),.clk(clk),.wout(w79_53));
	PE pe79_54(.x(x54),.w(w79_53),.acc(r79_53),.res(r79_54),.clk(clk),.wout(w79_54));
	PE pe79_55(.x(x55),.w(w79_54),.acc(r79_54),.res(r79_55),.clk(clk),.wout(w79_55));
	PE pe79_56(.x(x56),.w(w79_55),.acc(r79_55),.res(r79_56),.clk(clk),.wout(w79_56));
	PE pe79_57(.x(x57),.w(w79_56),.acc(r79_56),.res(r79_57),.clk(clk),.wout(w79_57));
	PE pe79_58(.x(x58),.w(w79_57),.acc(r79_57),.res(r79_58),.clk(clk),.wout(w79_58));
	PE pe79_59(.x(x59),.w(w79_58),.acc(r79_58),.res(r79_59),.clk(clk),.wout(w79_59));
	PE pe79_60(.x(x60),.w(w79_59),.acc(r79_59),.res(r79_60),.clk(clk),.wout(w79_60));
	PE pe79_61(.x(x61),.w(w79_60),.acc(r79_60),.res(r79_61),.clk(clk),.wout(w79_61));
	PE pe79_62(.x(x62),.w(w79_61),.acc(r79_61),.res(r79_62),.clk(clk),.wout(w79_62));
	PE pe79_63(.x(x63),.w(w79_62),.acc(r79_62),.res(r79_63),.clk(clk),.wout(w79_63));
	PE pe79_64(.x(x64),.w(w79_63),.acc(r79_63),.res(r79_64),.clk(clk),.wout(w79_64));
	PE pe79_65(.x(x65),.w(w79_64),.acc(r79_64),.res(r79_65),.clk(clk),.wout(w79_65));
	PE pe79_66(.x(x66),.w(w79_65),.acc(r79_65),.res(r79_66),.clk(clk),.wout(w79_66));
	PE pe79_67(.x(x67),.w(w79_66),.acc(r79_66),.res(r79_67),.clk(clk),.wout(w79_67));
	PE pe79_68(.x(x68),.w(w79_67),.acc(r79_67),.res(r79_68),.clk(clk),.wout(w79_68));
	PE pe79_69(.x(x69),.w(w79_68),.acc(r79_68),.res(r79_69),.clk(clk),.wout(w79_69));
	PE pe79_70(.x(x70),.w(w79_69),.acc(r79_69),.res(r79_70),.clk(clk),.wout(w79_70));
	PE pe79_71(.x(x71),.w(w79_70),.acc(r79_70),.res(r79_71),.clk(clk),.wout(w79_71));
	PE pe79_72(.x(x72),.w(w79_71),.acc(r79_71),.res(r79_72),.clk(clk),.wout(w79_72));
	PE pe79_73(.x(x73),.w(w79_72),.acc(r79_72),.res(r79_73),.clk(clk),.wout(w79_73));
	PE pe79_74(.x(x74),.w(w79_73),.acc(r79_73),.res(r79_74),.clk(clk),.wout(w79_74));
	PE pe79_75(.x(x75),.w(w79_74),.acc(r79_74),.res(r79_75),.clk(clk),.wout(w79_75));
	PE pe79_76(.x(x76),.w(w79_75),.acc(r79_75),.res(r79_76),.clk(clk),.wout(w79_76));
	PE pe79_77(.x(x77),.w(w79_76),.acc(r79_76),.res(r79_77),.clk(clk),.wout(w79_77));
	PE pe79_78(.x(x78),.w(w79_77),.acc(r79_77),.res(r79_78),.clk(clk),.wout(w79_78));
	PE pe79_79(.x(x79),.w(w79_78),.acc(r79_78),.res(r79_79),.clk(clk),.wout(w79_79));
	PE pe79_80(.x(x80),.w(w79_79),.acc(r79_79),.res(r79_80),.clk(clk),.wout(w79_80));
	PE pe79_81(.x(x81),.w(w79_80),.acc(r79_80),.res(r79_81),.clk(clk),.wout(w79_81));
	PE pe79_82(.x(x82),.w(w79_81),.acc(r79_81),.res(r79_82),.clk(clk),.wout(w79_82));
	PE pe79_83(.x(x83),.w(w79_82),.acc(r79_82),.res(r79_83),.clk(clk),.wout(w79_83));
	PE pe79_84(.x(x84),.w(w79_83),.acc(r79_83),.res(r79_84),.clk(clk),.wout(w79_84));
	PE pe79_85(.x(x85),.w(w79_84),.acc(r79_84),.res(r79_85),.clk(clk),.wout(w79_85));
	PE pe79_86(.x(x86),.w(w79_85),.acc(r79_85),.res(r79_86),.clk(clk),.wout(w79_86));
	PE pe79_87(.x(x87),.w(w79_86),.acc(r79_86),.res(r79_87),.clk(clk),.wout(w79_87));
	PE pe79_88(.x(x88),.w(w79_87),.acc(r79_87),.res(r79_88),.clk(clk),.wout(w79_88));
	PE pe79_89(.x(x89),.w(w79_88),.acc(r79_88),.res(r79_89),.clk(clk),.wout(w79_89));
	PE pe79_90(.x(x90),.w(w79_89),.acc(r79_89),.res(r79_90),.clk(clk),.wout(w79_90));
	PE pe79_91(.x(x91),.w(w79_90),.acc(r79_90),.res(r79_91),.clk(clk),.wout(w79_91));
	PE pe79_92(.x(x92),.w(w79_91),.acc(r79_91),.res(r79_92),.clk(clk),.wout(w79_92));
	PE pe79_93(.x(x93),.w(w79_92),.acc(r79_92),.res(r79_93),.clk(clk),.wout(w79_93));
	PE pe79_94(.x(x94),.w(w79_93),.acc(r79_93),.res(r79_94),.clk(clk),.wout(w79_94));
	PE pe79_95(.x(x95),.w(w79_94),.acc(r79_94),.res(r79_95),.clk(clk),.wout(w79_95));
	PE pe79_96(.x(x96),.w(w79_95),.acc(r79_95),.res(r79_96),.clk(clk),.wout(w79_96));
	PE pe79_97(.x(x97),.w(w79_96),.acc(r79_96),.res(r79_97),.clk(clk),.wout(w79_97));
	PE pe79_98(.x(x98),.w(w79_97),.acc(r79_97),.res(r79_98),.clk(clk),.wout(w79_98));
	PE pe79_99(.x(x99),.w(w79_98),.acc(r79_98),.res(r79_99),.clk(clk),.wout(w79_99));
	PE pe79_100(.x(x100),.w(w79_99),.acc(r79_99),.res(r79_100),.clk(clk),.wout(w79_100));
	PE pe79_101(.x(x101),.w(w79_100),.acc(r79_100),.res(r79_101),.clk(clk),.wout(w79_101));
	PE pe79_102(.x(x102),.w(w79_101),.acc(r79_101),.res(r79_102),.clk(clk),.wout(w79_102));
	PE pe79_103(.x(x103),.w(w79_102),.acc(r79_102),.res(r79_103),.clk(clk),.wout(w79_103));
	PE pe79_104(.x(x104),.w(w79_103),.acc(r79_103),.res(r79_104),.clk(clk),.wout(w79_104));
	PE pe79_105(.x(x105),.w(w79_104),.acc(r79_104),.res(r79_105),.clk(clk),.wout(w79_105));
	PE pe79_106(.x(x106),.w(w79_105),.acc(r79_105),.res(r79_106),.clk(clk),.wout(w79_106));
	PE pe79_107(.x(x107),.w(w79_106),.acc(r79_106),.res(r79_107),.clk(clk),.wout(w79_107));
	PE pe79_108(.x(x108),.w(w79_107),.acc(r79_107),.res(r79_108),.clk(clk),.wout(w79_108));
	PE pe79_109(.x(x109),.w(w79_108),.acc(r79_108),.res(r79_109),.clk(clk),.wout(w79_109));
	PE pe79_110(.x(x110),.w(w79_109),.acc(r79_109),.res(r79_110),.clk(clk),.wout(w79_110));
	PE pe79_111(.x(x111),.w(w79_110),.acc(r79_110),.res(r79_111),.clk(clk),.wout(w79_111));
	PE pe79_112(.x(x112),.w(w79_111),.acc(r79_111),.res(r79_112),.clk(clk),.wout(w79_112));
	PE pe79_113(.x(x113),.w(w79_112),.acc(r79_112),.res(r79_113),.clk(clk),.wout(w79_113));
	PE pe79_114(.x(x114),.w(w79_113),.acc(r79_113),.res(r79_114),.clk(clk),.wout(w79_114));
	PE pe79_115(.x(x115),.w(w79_114),.acc(r79_114),.res(r79_115),.clk(clk),.wout(w79_115));
	PE pe79_116(.x(x116),.w(w79_115),.acc(r79_115),.res(r79_116),.clk(clk),.wout(w79_116));
	PE pe79_117(.x(x117),.w(w79_116),.acc(r79_116),.res(r79_117),.clk(clk),.wout(w79_117));
	PE pe79_118(.x(x118),.w(w79_117),.acc(r79_117),.res(r79_118),.clk(clk),.wout(w79_118));
	PE pe79_119(.x(x119),.w(w79_118),.acc(r79_118),.res(r79_119),.clk(clk),.wout(w79_119));
	PE pe79_120(.x(x120),.w(w79_119),.acc(r79_119),.res(r79_120),.clk(clk),.wout(w79_120));
	PE pe79_121(.x(x121),.w(w79_120),.acc(r79_120),.res(r79_121),.clk(clk),.wout(w79_121));
	PE pe79_122(.x(x122),.w(w79_121),.acc(r79_121),.res(r79_122),.clk(clk),.wout(w79_122));
	PE pe79_123(.x(x123),.w(w79_122),.acc(r79_122),.res(r79_123),.clk(clk),.wout(w79_123));
	PE pe79_124(.x(x124),.w(w79_123),.acc(r79_123),.res(r79_124),.clk(clk),.wout(w79_124));
	PE pe79_125(.x(x125),.w(w79_124),.acc(r79_124),.res(r79_125),.clk(clk),.wout(w79_125));
	PE pe79_126(.x(x126),.w(w79_125),.acc(r79_125),.res(r79_126),.clk(clk),.wout(w79_126));
	PE pe79_127(.x(x127),.w(w79_126),.acc(r79_126),.res(result79),.clk(clk),.wout(weight79));

	PE pe80_0(.x(x0),.w(w80),.acc(32'h0),.res(r80_0),.clk(clk),.wout(w80_0));
	PE pe80_1(.x(x1),.w(w80_0),.acc(r80_0),.res(r80_1),.clk(clk),.wout(w80_1));
	PE pe80_2(.x(x2),.w(w80_1),.acc(r80_1),.res(r80_2),.clk(clk),.wout(w80_2));
	PE pe80_3(.x(x3),.w(w80_2),.acc(r80_2),.res(r80_3),.clk(clk),.wout(w80_3));
	PE pe80_4(.x(x4),.w(w80_3),.acc(r80_3),.res(r80_4),.clk(clk),.wout(w80_4));
	PE pe80_5(.x(x5),.w(w80_4),.acc(r80_4),.res(r80_5),.clk(clk),.wout(w80_5));
	PE pe80_6(.x(x6),.w(w80_5),.acc(r80_5),.res(r80_6),.clk(clk),.wout(w80_6));
	PE pe80_7(.x(x7),.w(w80_6),.acc(r80_6),.res(r80_7),.clk(clk),.wout(w80_7));
	PE pe80_8(.x(x8),.w(w80_7),.acc(r80_7),.res(r80_8),.clk(clk),.wout(w80_8));
	PE pe80_9(.x(x9),.w(w80_8),.acc(r80_8),.res(r80_9),.clk(clk),.wout(w80_9));
	PE pe80_10(.x(x10),.w(w80_9),.acc(r80_9),.res(r80_10),.clk(clk),.wout(w80_10));
	PE pe80_11(.x(x11),.w(w80_10),.acc(r80_10),.res(r80_11),.clk(clk),.wout(w80_11));
	PE pe80_12(.x(x12),.w(w80_11),.acc(r80_11),.res(r80_12),.clk(clk),.wout(w80_12));
	PE pe80_13(.x(x13),.w(w80_12),.acc(r80_12),.res(r80_13),.clk(clk),.wout(w80_13));
	PE pe80_14(.x(x14),.w(w80_13),.acc(r80_13),.res(r80_14),.clk(clk),.wout(w80_14));
	PE pe80_15(.x(x15),.w(w80_14),.acc(r80_14),.res(r80_15),.clk(clk),.wout(w80_15));
	PE pe80_16(.x(x16),.w(w80_15),.acc(r80_15),.res(r80_16),.clk(clk),.wout(w80_16));
	PE pe80_17(.x(x17),.w(w80_16),.acc(r80_16),.res(r80_17),.clk(clk),.wout(w80_17));
	PE pe80_18(.x(x18),.w(w80_17),.acc(r80_17),.res(r80_18),.clk(clk),.wout(w80_18));
	PE pe80_19(.x(x19),.w(w80_18),.acc(r80_18),.res(r80_19),.clk(clk),.wout(w80_19));
	PE pe80_20(.x(x20),.w(w80_19),.acc(r80_19),.res(r80_20),.clk(clk),.wout(w80_20));
	PE pe80_21(.x(x21),.w(w80_20),.acc(r80_20),.res(r80_21),.clk(clk),.wout(w80_21));
	PE pe80_22(.x(x22),.w(w80_21),.acc(r80_21),.res(r80_22),.clk(clk),.wout(w80_22));
	PE pe80_23(.x(x23),.w(w80_22),.acc(r80_22),.res(r80_23),.clk(clk),.wout(w80_23));
	PE pe80_24(.x(x24),.w(w80_23),.acc(r80_23),.res(r80_24),.clk(clk),.wout(w80_24));
	PE pe80_25(.x(x25),.w(w80_24),.acc(r80_24),.res(r80_25),.clk(clk),.wout(w80_25));
	PE pe80_26(.x(x26),.w(w80_25),.acc(r80_25),.res(r80_26),.clk(clk),.wout(w80_26));
	PE pe80_27(.x(x27),.w(w80_26),.acc(r80_26),.res(r80_27),.clk(clk),.wout(w80_27));
	PE pe80_28(.x(x28),.w(w80_27),.acc(r80_27),.res(r80_28),.clk(clk),.wout(w80_28));
	PE pe80_29(.x(x29),.w(w80_28),.acc(r80_28),.res(r80_29),.clk(clk),.wout(w80_29));
	PE pe80_30(.x(x30),.w(w80_29),.acc(r80_29),.res(r80_30),.clk(clk),.wout(w80_30));
	PE pe80_31(.x(x31),.w(w80_30),.acc(r80_30),.res(r80_31),.clk(clk),.wout(w80_31));
	PE pe80_32(.x(x32),.w(w80_31),.acc(r80_31),.res(r80_32),.clk(clk),.wout(w80_32));
	PE pe80_33(.x(x33),.w(w80_32),.acc(r80_32),.res(r80_33),.clk(clk),.wout(w80_33));
	PE pe80_34(.x(x34),.w(w80_33),.acc(r80_33),.res(r80_34),.clk(clk),.wout(w80_34));
	PE pe80_35(.x(x35),.w(w80_34),.acc(r80_34),.res(r80_35),.clk(clk),.wout(w80_35));
	PE pe80_36(.x(x36),.w(w80_35),.acc(r80_35),.res(r80_36),.clk(clk),.wout(w80_36));
	PE pe80_37(.x(x37),.w(w80_36),.acc(r80_36),.res(r80_37),.clk(clk),.wout(w80_37));
	PE pe80_38(.x(x38),.w(w80_37),.acc(r80_37),.res(r80_38),.clk(clk),.wout(w80_38));
	PE pe80_39(.x(x39),.w(w80_38),.acc(r80_38),.res(r80_39),.clk(clk),.wout(w80_39));
	PE pe80_40(.x(x40),.w(w80_39),.acc(r80_39),.res(r80_40),.clk(clk),.wout(w80_40));
	PE pe80_41(.x(x41),.w(w80_40),.acc(r80_40),.res(r80_41),.clk(clk),.wout(w80_41));
	PE pe80_42(.x(x42),.w(w80_41),.acc(r80_41),.res(r80_42),.clk(clk),.wout(w80_42));
	PE pe80_43(.x(x43),.w(w80_42),.acc(r80_42),.res(r80_43),.clk(clk),.wout(w80_43));
	PE pe80_44(.x(x44),.w(w80_43),.acc(r80_43),.res(r80_44),.clk(clk),.wout(w80_44));
	PE pe80_45(.x(x45),.w(w80_44),.acc(r80_44),.res(r80_45),.clk(clk),.wout(w80_45));
	PE pe80_46(.x(x46),.w(w80_45),.acc(r80_45),.res(r80_46),.clk(clk),.wout(w80_46));
	PE pe80_47(.x(x47),.w(w80_46),.acc(r80_46),.res(r80_47),.clk(clk),.wout(w80_47));
	PE pe80_48(.x(x48),.w(w80_47),.acc(r80_47),.res(r80_48),.clk(clk),.wout(w80_48));
	PE pe80_49(.x(x49),.w(w80_48),.acc(r80_48),.res(r80_49),.clk(clk),.wout(w80_49));
	PE pe80_50(.x(x50),.w(w80_49),.acc(r80_49),.res(r80_50),.clk(clk),.wout(w80_50));
	PE pe80_51(.x(x51),.w(w80_50),.acc(r80_50),.res(r80_51),.clk(clk),.wout(w80_51));
	PE pe80_52(.x(x52),.w(w80_51),.acc(r80_51),.res(r80_52),.clk(clk),.wout(w80_52));
	PE pe80_53(.x(x53),.w(w80_52),.acc(r80_52),.res(r80_53),.clk(clk),.wout(w80_53));
	PE pe80_54(.x(x54),.w(w80_53),.acc(r80_53),.res(r80_54),.clk(clk),.wout(w80_54));
	PE pe80_55(.x(x55),.w(w80_54),.acc(r80_54),.res(r80_55),.clk(clk),.wout(w80_55));
	PE pe80_56(.x(x56),.w(w80_55),.acc(r80_55),.res(r80_56),.clk(clk),.wout(w80_56));
	PE pe80_57(.x(x57),.w(w80_56),.acc(r80_56),.res(r80_57),.clk(clk),.wout(w80_57));
	PE pe80_58(.x(x58),.w(w80_57),.acc(r80_57),.res(r80_58),.clk(clk),.wout(w80_58));
	PE pe80_59(.x(x59),.w(w80_58),.acc(r80_58),.res(r80_59),.clk(clk),.wout(w80_59));
	PE pe80_60(.x(x60),.w(w80_59),.acc(r80_59),.res(r80_60),.clk(clk),.wout(w80_60));
	PE pe80_61(.x(x61),.w(w80_60),.acc(r80_60),.res(r80_61),.clk(clk),.wout(w80_61));
	PE pe80_62(.x(x62),.w(w80_61),.acc(r80_61),.res(r80_62),.clk(clk),.wout(w80_62));
	PE pe80_63(.x(x63),.w(w80_62),.acc(r80_62),.res(r80_63),.clk(clk),.wout(w80_63));
	PE pe80_64(.x(x64),.w(w80_63),.acc(r80_63),.res(r80_64),.clk(clk),.wout(w80_64));
	PE pe80_65(.x(x65),.w(w80_64),.acc(r80_64),.res(r80_65),.clk(clk),.wout(w80_65));
	PE pe80_66(.x(x66),.w(w80_65),.acc(r80_65),.res(r80_66),.clk(clk),.wout(w80_66));
	PE pe80_67(.x(x67),.w(w80_66),.acc(r80_66),.res(r80_67),.clk(clk),.wout(w80_67));
	PE pe80_68(.x(x68),.w(w80_67),.acc(r80_67),.res(r80_68),.clk(clk),.wout(w80_68));
	PE pe80_69(.x(x69),.w(w80_68),.acc(r80_68),.res(r80_69),.clk(clk),.wout(w80_69));
	PE pe80_70(.x(x70),.w(w80_69),.acc(r80_69),.res(r80_70),.clk(clk),.wout(w80_70));
	PE pe80_71(.x(x71),.w(w80_70),.acc(r80_70),.res(r80_71),.clk(clk),.wout(w80_71));
	PE pe80_72(.x(x72),.w(w80_71),.acc(r80_71),.res(r80_72),.clk(clk),.wout(w80_72));
	PE pe80_73(.x(x73),.w(w80_72),.acc(r80_72),.res(r80_73),.clk(clk),.wout(w80_73));
	PE pe80_74(.x(x74),.w(w80_73),.acc(r80_73),.res(r80_74),.clk(clk),.wout(w80_74));
	PE pe80_75(.x(x75),.w(w80_74),.acc(r80_74),.res(r80_75),.clk(clk),.wout(w80_75));
	PE pe80_76(.x(x76),.w(w80_75),.acc(r80_75),.res(r80_76),.clk(clk),.wout(w80_76));
	PE pe80_77(.x(x77),.w(w80_76),.acc(r80_76),.res(r80_77),.clk(clk),.wout(w80_77));
	PE pe80_78(.x(x78),.w(w80_77),.acc(r80_77),.res(r80_78),.clk(clk),.wout(w80_78));
	PE pe80_79(.x(x79),.w(w80_78),.acc(r80_78),.res(r80_79),.clk(clk),.wout(w80_79));
	PE pe80_80(.x(x80),.w(w80_79),.acc(r80_79),.res(r80_80),.clk(clk),.wout(w80_80));
	PE pe80_81(.x(x81),.w(w80_80),.acc(r80_80),.res(r80_81),.clk(clk),.wout(w80_81));
	PE pe80_82(.x(x82),.w(w80_81),.acc(r80_81),.res(r80_82),.clk(clk),.wout(w80_82));
	PE pe80_83(.x(x83),.w(w80_82),.acc(r80_82),.res(r80_83),.clk(clk),.wout(w80_83));
	PE pe80_84(.x(x84),.w(w80_83),.acc(r80_83),.res(r80_84),.clk(clk),.wout(w80_84));
	PE pe80_85(.x(x85),.w(w80_84),.acc(r80_84),.res(r80_85),.clk(clk),.wout(w80_85));
	PE pe80_86(.x(x86),.w(w80_85),.acc(r80_85),.res(r80_86),.clk(clk),.wout(w80_86));
	PE pe80_87(.x(x87),.w(w80_86),.acc(r80_86),.res(r80_87),.clk(clk),.wout(w80_87));
	PE pe80_88(.x(x88),.w(w80_87),.acc(r80_87),.res(r80_88),.clk(clk),.wout(w80_88));
	PE pe80_89(.x(x89),.w(w80_88),.acc(r80_88),.res(r80_89),.clk(clk),.wout(w80_89));
	PE pe80_90(.x(x90),.w(w80_89),.acc(r80_89),.res(r80_90),.clk(clk),.wout(w80_90));
	PE pe80_91(.x(x91),.w(w80_90),.acc(r80_90),.res(r80_91),.clk(clk),.wout(w80_91));
	PE pe80_92(.x(x92),.w(w80_91),.acc(r80_91),.res(r80_92),.clk(clk),.wout(w80_92));
	PE pe80_93(.x(x93),.w(w80_92),.acc(r80_92),.res(r80_93),.clk(clk),.wout(w80_93));
	PE pe80_94(.x(x94),.w(w80_93),.acc(r80_93),.res(r80_94),.clk(clk),.wout(w80_94));
	PE pe80_95(.x(x95),.w(w80_94),.acc(r80_94),.res(r80_95),.clk(clk),.wout(w80_95));
	PE pe80_96(.x(x96),.w(w80_95),.acc(r80_95),.res(r80_96),.clk(clk),.wout(w80_96));
	PE pe80_97(.x(x97),.w(w80_96),.acc(r80_96),.res(r80_97),.clk(clk),.wout(w80_97));
	PE pe80_98(.x(x98),.w(w80_97),.acc(r80_97),.res(r80_98),.clk(clk),.wout(w80_98));
	PE pe80_99(.x(x99),.w(w80_98),.acc(r80_98),.res(r80_99),.clk(clk),.wout(w80_99));
	PE pe80_100(.x(x100),.w(w80_99),.acc(r80_99),.res(r80_100),.clk(clk),.wout(w80_100));
	PE pe80_101(.x(x101),.w(w80_100),.acc(r80_100),.res(r80_101),.clk(clk),.wout(w80_101));
	PE pe80_102(.x(x102),.w(w80_101),.acc(r80_101),.res(r80_102),.clk(clk),.wout(w80_102));
	PE pe80_103(.x(x103),.w(w80_102),.acc(r80_102),.res(r80_103),.clk(clk),.wout(w80_103));
	PE pe80_104(.x(x104),.w(w80_103),.acc(r80_103),.res(r80_104),.clk(clk),.wout(w80_104));
	PE pe80_105(.x(x105),.w(w80_104),.acc(r80_104),.res(r80_105),.clk(clk),.wout(w80_105));
	PE pe80_106(.x(x106),.w(w80_105),.acc(r80_105),.res(r80_106),.clk(clk),.wout(w80_106));
	PE pe80_107(.x(x107),.w(w80_106),.acc(r80_106),.res(r80_107),.clk(clk),.wout(w80_107));
	PE pe80_108(.x(x108),.w(w80_107),.acc(r80_107),.res(r80_108),.clk(clk),.wout(w80_108));
	PE pe80_109(.x(x109),.w(w80_108),.acc(r80_108),.res(r80_109),.clk(clk),.wout(w80_109));
	PE pe80_110(.x(x110),.w(w80_109),.acc(r80_109),.res(r80_110),.clk(clk),.wout(w80_110));
	PE pe80_111(.x(x111),.w(w80_110),.acc(r80_110),.res(r80_111),.clk(clk),.wout(w80_111));
	PE pe80_112(.x(x112),.w(w80_111),.acc(r80_111),.res(r80_112),.clk(clk),.wout(w80_112));
	PE pe80_113(.x(x113),.w(w80_112),.acc(r80_112),.res(r80_113),.clk(clk),.wout(w80_113));
	PE pe80_114(.x(x114),.w(w80_113),.acc(r80_113),.res(r80_114),.clk(clk),.wout(w80_114));
	PE pe80_115(.x(x115),.w(w80_114),.acc(r80_114),.res(r80_115),.clk(clk),.wout(w80_115));
	PE pe80_116(.x(x116),.w(w80_115),.acc(r80_115),.res(r80_116),.clk(clk),.wout(w80_116));
	PE pe80_117(.x(x117),.w(w80_116),.acc(r80_116),.res(r80_117),.clk(clk),.wout(w80_117));
	PE pe80_118(.x(x118),.w(w80_117),.acc(r80_117),.res(r80_118),.clk(clk),.wout(w80_118));
	PE pe80_119(.x(x119),.w(w80_118),.acc(r80_118),.res(r80_119),.clk(clk),.wout(w80_119));
	PE pe80_120(.x(x120),.w(w80_119),.acc(r80_119),.res(r80_120),.clk(clk),.wout(w80_120));
	PE pe80_121(.x(x121),.w(w80_120),.acc(r80_120),.res(r80_121),.clk(clk),.wout(w80_121));
	PE pe80_122(.x(x122),.w(w80_121),.acc(r80_121),.res(r80_122),.clk(clk),.wout(w80_122));
	PE pe80_123(.x(x123),.w(w80_122),.acc(r80_122),.res(r80_123),.clk(clk),.wout(w80_123));
	PE pe80_124(.x(x124),.w(w80_123),.acc(r80_123),.res(r80_124),.clk(clk),.wout(w80_124));
	PE pe80_125(.x(x125),.w(w80_124),.acc(r80_124),.res(r80_125),.clk(clk),.wout(w80_125));
	PE pe80_126(.x(x126),.w(w80_125),.acc(r80_125),.res(r80_126),.clk(clk),.wout(w80_126));
	PE pe80_127(.x(x127),.w(w80_126),.acc(r80_126),.res(result80),.clk(clk),.wout(weight80));

	PE pe81_0(.x(x0),.w(w81),.acc(32'h0),.res(r81_0),.clk(clk),.wout(w81_0));
	PE pe81_1(.x(x1),.w(w81_0),.acc(r81_0),.res(r81_1),.clk(clk),.wout(w81_1));
	PE pe81_2(.x(x2),.w(w81_1),.acc(r81_1),.res(r81_2),.clk(clk),.wout(w81_2));
	PE pe81_3(.x(x3),.w(w81_2),.acc(r81_2),.res(r81_3),.clk(clk),.wout(w81_3));
	PE pe81_4(.x(x4),.w(w81_3),.acc(r81_3),.res(r81_4),.clk(clk),.wout(w81_4));
	PE pe81_5(.x(x5),.w(w81_4),.acc(r81_4),.res(r81_5),.clk(clk),.wout(w81_5));
	PE pe81_6(.x(x6),.w(w81_5),.acc(r81_5),.res(r81_6),.clk(clk),.wout(w81_6));
	PE pe81_7(.x(x7),.w(w81_6),.acc(r81_6),.res(r81_7),.clk(clk),.wout(w81_7));
	PE pe81_8(.x(x8),.w(w81_7),.acc(r81_7),.res(r81_8),.clk(clk),.wout(w81_8));
	PE pe81_9(.x(x9),.w(w81_8),.acc(r81_8),.res(r81_9),.clk(clk),.wout(w81_9));
	PE pe81_10(.x(x10),.w(w81_9),.acc(r81_9),.res(r81_10),.clk(clk),.wout(w81_10));
	PE pe81_11(.x(x11),.w(w81_10),.acc(r81_10),.res(r81_11),.clk(clk),.wout(w81_11));
	PE pe81_12(.x(x12),.w(w81_11),.acc(r81_11),.res(r81_12),.clk(clk),.wout(w81_12));
	PE pe81_13(.x(x13),.w(w81_12),.acc(r81_12),.res(r81_13),.clk(clk),.wout(w81_13));
	PE pe81_14(.x(x14),.w(w81_13),.acc(r81_13),.res(r81_14),.clk(clk),.wout(w81_14));
	PE pe81_15(.x(x15),.w(w81_14),.acc(r81_14),.res(r81_15),.clk(clk),.wout(w81_15));
	PE pe81_16(.x(x16),.w(w81_15),.acc(r81_15),.res(r81_16),.clk(clk),.wout(w81_16));
	PE pe81_17(.x(x17),.w(w81_16),.acc(r81_16),.res(r81_17),.clk(clk),.wout(w81_17));
	PE pe81_18(.x(x18),.w(w81_17),.acc(r81_17),.res(r81_18),.clk(clk),.wout(w81_18));
	PE pe81_19(.x(x19),.w(w81_18),.acc(r81_18),.res(r81_19),.clk(clk),.wout(w81_19));
	PE pe81_20(.x(x20),.w(w81_19),.acc(r81_19),.res(r81_20),.clk(clk),.wout(w81_20));
	PE pe81_21(.x(x21),.w(w81_20),.acc(r81_20),.res(r81_21),.clk(clk),.wout(w81_21));
	PE pe81_22(.x(x22),.w(w81_21),.acc(r81_21),.res(r81_22),.clk(clk),.wout(w81_22));
	PE pe81_23(.x(x23),.w(w81_22),.acc(r81_22),.res(r81_23),.clk(clk),.wout(w81_23));
	PE pe81_24(.x(x24),.w(w81_23),.acc(r81_23),.res(r81_24),.clk(clk),.wout(w81_24));
	PE pe81_25(.x(x25),.w(w81_24),.acc(r81_24),.res(r81_25),.clk(clk),.wout(w81_25));
	PE pe81_26(.x(x26),.w(w81_25),.acc(r81_25),.res(r81_26),.clk(clk),.wout(w81_26));
	PE pe81_27(.x(x27),.w(w81_26),.acc(r81_26),.res(r81_27),.clk(clk),.wout(w81_27));
	PE pe81_28(.x(x28),.w(w81_27),.acc(r81_27),.res(r81_28),.clk(clk),.wout(w81_28));
	PE pe81_29(.x(x29),.w(w81_28),.acc(r81_28),.res(r81_29),.clk(clk),.wout(w81_29));
	PE pe81_30(.x(x30),.w(w81_29),.acc(r81_29),.res(r81_30),.clk(clk),.wout(w81_30));
	PE pe81_31(.x(x31),.w(w81_30),.acc(r81_30),.res(r81_31),.clk(clk),.wout(w81_31));
	PE pe81_32(.x(x32),.w(w81_31),.acc(r81_31),.res(r81_32),.clk(clk),.wout(w81_32));
	PE pe81_33(.x(x33),.w(w81_32),.acc(r81_32),.res(r81_33),.clk(clk),.wout(w81_33));
	PE pe81_34(.x(x34),.w(w81_33),.acc(r81_33),.res(r81_34),.clk(clk),.wout(w81_34));
	PE pe81_35(.x(x35),.w(w81_34),.acc(r81_34),.res(r81_35),.clk(clk),.wout(w81_35));
	PE pe81_36(.x(x36),.w(w81_35),.acc(r81_35),.res(r81_36),.clk(clk),.wout(w81_36));
	PE pe81_37(.x(x37),.w(w81_36),.acc(r81_36),.res(r81_37),.clk(clk),.wout(w81_37));
	PE pe81_38(.x(x38),.w(w81_37),.acc(r81_37),.res(r81_38),.clk(clk),.wout(w81_38));
	PE pe81_39(.x(x39),.w(w81_38),.acc(r81_38),.res(r81_39),.clk(clk),.wout(w81_39));
	PE pe81_40(.x(x40),.w(w81_39),.acc(r81_39),.res(r81_40),.clk(clk),.wout(w81_40));
	PE pe81_41(.x(x41),.w(w81_40),.acc(r81_40),.res(r81_41),.clk(clk),.wout(w81_41));
	PE pe81_42(.x(x42),.w(w81_41),.acc(r81_41),.res(r81_42),.clk(clk),.wout(w81_42));
	PE pe81_43(.x(x43),.w(w81_42),.acc(r81_42),.res(r81_43),.clk(clk),.wout(w81_43));
	PE pe81_44(.x(x44),.w(w81_43),.acc(r81_43),.res(r81_44),.clk(clk),.wout(w81_44));
	PE pe81_45(.x(x45),.w(w81_44),.acc(r81_44),.res(r81_45),.clk(clk),.wout(w81_45));
	PE pe81_46(.x(x46),.w(w81_45),.acc(r81_45),.res(r81_46),.clk(clk),.wout(w81_46));
	PE pe81_47(.x(x47),.w(w81_46),.acc(r81_46),.res(r81_47),.clk(clk),.wout(w81_47));
	PE pe81_48(.x(x48),.w(w81_47),.acc(r81_47),.res(r81_48),.clk(clk),.wout(w81_48));
	PE pe81_49(.x(x49),.w(w81_48),.acc(r81_48),.res(r81_49),.clk(clk),.wout(w81_49));
	PE pe81_50(.x(x50),.w(w81_49),.acc(r81_49),.res(r81_50),.clk(clk),.wout(w81_50));
	PE pe81_51(.x(x51),.w(w81_50),.acc(r81_50),.res(r81_51),.clk(clk),.wout(w81_51));
	PE pe81_52(.x(x52),.w(w81_51),.acc(r81_51),.res(r81_52),.clk(clk),.wout(w81_52));
	PE pe81_53(.x(x53),.w(w81_52),.acc(r81_52),.res(r81_53),.clk(clk),.wout(w81_53));
	PE pe81_54(.x(x54),.w(w81_53),.acc(r81_53),.res(r81_54),.clk(clk),.wout(w81_54));
	PE pe81_55(.x(x55),.w(w81_54),.acc(r81_54),.res(r81_55),.clk(clk),.wout(w81_55));
	PE pe81_56(.x(x56),.w(w81_55),.acc(r81_55),.res(r81_56),.clk(clk),.wout(w81_56));
	PE pe81_57(.x(x57),.w(w81_56),.acc(r81_56),.res(r81_57),.clk(clk),.wout(w81_57));
	PE pe81_58(.x(x58),.w(w81_57),.acc(r81_57),.res(r81_58),.clk(clk),.wout(w81_58));
	PE pe81_59(.x(x59),.w(w81_58),.acc(r81_58),.res(r81_59),.clk(clk),.wout(w81_59));
	PE pe81_60(.x(x60),.w(w81_59),.acc(r81_59),.res(r81_60),.clk(clk),.wout(w81_60));
	PE pe81_61(.x(x61),.w(w81_60),.acc(r81_60),.res(r81_61),.clk(clk),.wout(w81_61));
	PE pe81_62(.x(x62),.w(w81_61),.acc(r81_61),.res(r81_62),.clk(clk),.wout(w81_62));
	PE pe81_63(.x(x63),.w(w81_62),.acc(r81_62),.res(r81_63),.clk(clk),.wout(w81_63));
	PE pe81_64(.x(x64),.w(w81_63),.acc(r81_63),.res(r81_64),.clk(clk),.wout(w81_64));
	PE pe81_65(.x(x65),.w(w81_64),.acc(r81_64),.res(r81_65),.clk(clk),.wout(w81_65));
	PE pe81_66(.x(x66),.w(w81_65),.acc(r81_65),.res(r81_66),.clk(clk),.wout(w81_66));
	PE pe81_67(.x(x67),.w(w81_66),.acc(r81_66),.res(r81_67),.clk(clk),.wout(w81_67));
	PE pe81_68(.x(x68),.w(w81_67),.acc(r81_67),.res(r81_68),.clk(clk),.wout(w81_68));
	PE pe81_69(.x(x69),.w(w81_68),.acc(r81_68),.res(r81_69),.clk(clk),.wout(w81_69));
	PE pe81_70(.x(x70),.w(w81_69),.acc(r81_69),.res(r81_70),.clk(clk),.wout(w81_70));
	PE pe81_71(.x(x71),.w(w81_70),.acc(r81_70),.res(r81_71),.clk(clk),.wout(w81_71));
	PE pe81_72(.x(x72),.w(w81_71),.acc(r81_71),.res(r81_72),.clk(clk),.wout(w81_72));
	PE pe81_73(.x(x73),.w(w81_72),.acc(r81_72),.res(r81_73),.clk(clk),.wout(w81_73));
	PE pe81_74(.x(x74),.w(w81_73),.acc(r81_73),.res(r81_74),.clk(clk),.wout(w81_74));
	PE pe81_75(.x(x75),.w(w81_74),.acc(r81_74),.res(r81_75),.clk(clk),.wout(w81_75));
	PE pe81_76(.x(x76),.w(w81_75),.acc(r81_75),.res(r81_76),.clk(clk),.wout(w81_76));
	PE pe81_77(.x(x77),.w(w81_76),.acc(r81_76),.res(r81_77),.clk(clk),.wout(w81_77));
	PE pe81_78(.x(x78),.w(w81_77),.acc(r81_77),.res(r81_78),.clk(clk),.wout(w81_78));
	PE pe81_79(.x(x79),.w(w81_78),.acc(r81_78),.res(r81_79),.clk(clk),.wout(w81_79));
	PE pe81_80(.x(x80),.w(w81_79),.acc(r81_79),.res(r81_80),.clk(clk),.wout(w81_80));
	PE pe81_81(.x(x81),.w(w81_80),.acc(r81_80),.res(r81_81),.clk(clk),.wout(w81_81));
	PE pe81_82(.x(x82),.w(w81_81),.acc(r81_81),.res(r81_82),.clk(clk),.wout(w81_82));
	PE pe81_83(.x(x83),.w(w81_82),.acc(r81_82),.res(r81_83),.clk(clk),.wout(w81_83));
	PE pe81_84(.x(x84),.w(w81_83),.acc(r81_83),.res(r81_84),.clk(clk),.wout(w81_84));
	PE pe81_85(.x(x85),.w(w81_84),.acc(r81_84),.res(r81_85),.clk(clk),.wout(w81_85));
	PE pe81_86(.x(x86),.w(w81_85),.acc(r81_85),.res(r81_86),.clk(clk),.wout(w81_86));
	PE pe81_87(.x(x87),.w(w81_86),.acc(r81_86),.res(r81_87),.clk(clk),.wout(w81_87));
	PE pe81_88(.x(x88),.w(w81_87),.acc(r81_87),.res(r81_88),.clk(clk),.wout(w81_88));
	PE pe81_89(.x(x89),.w(w81_88),.acc(r81_88),.res(r81_89),.clk(clk),.wout(w81_89));
	PE pe81_90(.x(x90),.w(w81_89),.acc(r81_89),.res(r81_90),.clk(clk),.wout(w81_90));
	PE pe81_91(.x(x91),.w(w81_90),.acc(r81_90),.res(r81_91),.clk(clk),.wout(w81_91));
	PE pe81_92(.x(x92),.w(w81_91),.acc(r81_91),.res(r81_92),.clk(clk),.wout(w81_92));
	PE pe81_93(.x(x93),.w(w81_92),.acc(r81_92),.res(r81_93),.clk(clk),.wout(w81_93));
	PE pe81_94(.x(x94),.w(w81_93),.acc(r81_93),.res(r81_94),.clk(clk),.wout(w81_94));
	PE pe81_95(.x(x95),.w(w81_94),.acc(r81_94),.res(r81_95),.clk(clk),.wout(w81_95));
	PE pe81_96(.x(x96),.w(w81_95),.acc(r81_95),.res(r81_96),.clk(clk),.wout(w81_96));
	PE pe81_97(.x(x97),.w(w81_96),.acc(r81_96),.res(r81_97),.clk(clk),.wout(w81_97));
	PE pe81_98(.x(x98),.w(w81_97),.acc(r81_97),.res(r81_98),.clk(clk),.wout(w81_98));
	PE pe81_99(.x(x99),.w(w81_98),.acc(r81_98),.res(r81_99),.clk(clk),.wout(w81_99));
	PE pe81_100(.x(x100),.w(w81_99),.acc(r81_99),.res(r81_100),.clk(clk),.wout(w81_100));
	PE pe81_101(.x(x101),.w(w81_100),.acc(r81_100),.res(r81_101),.clk(clk),.wout(w81_101));
	PE pe81_102(.x(x102),.w(w81_101),.acc(r81_101),.res(r81_102),.clk(clk),.wout(w81_102));
	PE pe81_103(.x(x103),.w(w81_102),.acc(r81_102),.res(r81_103),.clk(clk),.wout(w81_103));
	PE pe81_104(.x(x104),.w(w81_103),.acc(r81_103),.res(r81_104),.clk(clk),.wout(w81_104));
	PE pe81_105(.x(x105),.w(w81_104),.acc(r81_104),.res(r81_105),.clk(clk),.wout(w81_105));
	PE pe81_106(.x(x106),.w(w81_105),.acc(r81_105),.res(r81_106),.clk(clk),.wout(w81_106));
	PE pe81_107(.x(x107),.w(w81_106),.acc(r81_106),.res(r81_107),.clk(clk),.wout(w81_107));
	PE pe81_108(.x(x108),.w(w81_107),.acc(r81_107),.res(r81_108),.clk(clk),.wout(w81_108));
	PE pe81_109(.x(x109),.w(w81_108),.acc(r81_108),.res(r81_109),.clk(clk),.wout(w81_109));
	PE pe81_110(.x(x110),.w(w81_109),.acc(r81_109),.res(r81_110),.clk(clk),.wout(w81_110));
	PE pe81_111(.x(x111),.w(w81_110),.acc(r81_110),.res(r81_111),.clk(clk),.wout(w81_111));
	PE pe81_112(.x(x112),.w(w81_111),.acc(r81_111),.res(r81_112),.clk(clk),.wout(w81_112));
	PE pe81_113(.x(x113),.w(w81_112),.acc(r81_112),.res(r81_113),.clk(clk),.wout(w81_113));
	PE pe81_114(.x(x114),.w(w81_113),.acc(r81_113),.res(r81_114),.clk(clk),.wout(w81_114));
	PE pe81_115(.x(x115),.w(w81_114),.acc(r81_114),.res(r81_115),.clk(clk),.wout(w81_115));
	PE pe81_116(.x(x116),.w(w81_115),.acc(r81_115),.res(r81_116),.clk(clk),.wout(w81_116));
	PE pe81_117(.x(x117),.w(w81_116),.acc(r81_116),.res(r81_117),.clk(clk),.wout(w81_117));
	PE pe81_118(.x(x118),.w(w81_117),.acc(r81_117),.res(r81_118),.clk(clk),.wout(w81_118));
	PE pe81_119(.x(x119),.w(w81_118),.acc(r81_118),.res(r81_119),.clk(clk),.wout(w81_119));
	PE pe81_120(.x(x120),.w(w81_119),.acc(r81_119),.res(r81_120),.clk(clk),.wout(w81_120));
	PE pe81_121(.x(x121),.w(w81_120),.acc(r81_120),.res(r81_121),.clk(clk),.wout(w81_121));
	PE pe81_122(.x(x122),.w(w81_121),.acc(r81_121),.res(r81_122),.clk(clk),.wout(w81_122));
	PE pe81_123(.x(x123),.w(w81_122),.acc(r81_122),.res(r81_123),.clk(clk),.wout(w81_123));
	PE pe81_124(.x(x124),.w(w81_123),.acc(r81_123),.res(r81_124),.clk(clk),.wout(w81_124));
	PE pe81_125(.x(x125),.w(w81_124),.acc(r81_124),.res(r81_125),.clk(clk),.wout(w81_125));
	PE pe81_126(.x(x126),.w(w81_125),.acc(r81_125),.res(r81_126),.clk(clk),.wout(w81_126));
	PE pe81_127(.x(x127),.w(w81_126),.acc(r81_126),.res(result81),.clk(clk),.wout(weight81));

	PE pe82_0(.x(x0),.w(w82),.acc(32'h0),.res(r82_0),.clk(clk),.wout(w82_0));
	PE pe82_1(.x(x1),.w(w82_0),.acc(r82_0),.res(r82_1),.clk(clk),.wout(w82_1));
	PE pe82_2(.x(x2),.w(w82_1),.acc(r82_1),.res(r82_2),.clk(clk),.wout(w82_2));
	PE pe82_3(.x(x3),.w(w82_2),.acc(r82_2),.res(r82_3),.clk(clk),.wout(w82_3));
	PE pe82_4(.x(x4),.w(w82_3),.acc(r82_3),.res(r82_4),.clk(clk),.wout(w82_4));
	PE pe82_5(.x(x5),.w(w82_4),.acc(r82_4),.res(r82_5),.clk(clk),.wout(w82_5));
	PE pe82_6(.x(x6),.w(w82_5),.acc(r82_5),.res(r82_6),.clk(clk),.wout(w82_6));
	PE pe82_7(.x(x7),.w(w82_6),.acc(r82_6),.res(r82_7),.clk(clk),.wout(w82_7));
	PE pe82_8(.x(x8),.w(w82_7),.acc(r82_7),.res(r82_8),.clk(clk),.wout(w82_8));
	PE pe82_9(.x(x9),.w(w82_8),.acc(r82_8),.res(r82_9),.clk(clk),.wout(w82_9));
	PE pe82_10(.x(x10),.w(w82_9),.acc(r82_9),.res(r82_10),.clk(clk),.wout(w82_10));
	PE pe82_11(.x(x11),.w(w82_10),.acc(r82_10),.res(r82_11),.clk(clk),.wout(w82_11));
	PE pe82_12(.x(x12),.w(w82_11),.acc(r82_11),.res(r82_12),.clk(clk),.wout(w82_12));
	PE pe82_13(.x(x13),.w(w82_12),.acc(r82_12),.res(r82_13),.clk(clk),.wout(w82_13));
	PE pe82_14(.x(x14),.w(w82_13),.acc(r82_13),.res(r82_14),.clk(clk),.wout(w82_14));
	PE pe82_15(.x(x15),.w(w82_14),.acc(r82_14),.res(r82_15),.clk(clk),.wout(w82_15));
	PE pe82_16(.x(x16),.w(w82_15),.acc(r82_15),.res(r82_16),.clk(clk),.wout(w82_16));
	PE pe82_17(.x(x17),.w(w82_16),.acc(r82_16),.res(r82_17),.clk(clk),.wout(w82_17));
	PE pe82_18(.x(x18),.w(w82_17),.acc(r82_17),.res(r82_18),.clk(clk),.wout(w82_18));
	PE pe82_19(.x(x19),.w(w82_18),.acc(r82_18),.res(r82_19),.clk(clk),.wout(w82_19));
	PE pe82_20(.x(x20),.w(w82_19),.acc(r82_19),.res(r82_20),.clk(clk),.wout(w82_20));
	PE pe82_21(.x(x21),.w(w82_20),.acc(r82_20),.res(r82_21),.clk(clk),.wout(w82_21));
	PE pe82_22(.x(x22),.w(w82_21),.acc(r82_21),.res(r82_22),.clk(clk),.wout(w82_22));
	PE pe82_23(.x(x23),.w(w82_22),.acc(r82_22),.res(r82_23),.clk(clk),.wout(w82_23));
	PE pe82_24(.x(x24),.w(w82_23),.acc(r82_23),.res(r82_24),.clk(clk),.wout(w82_24));
	PE pe82_25(.x(x25),.w(w82_24),.acc(r82_24),.res(r82_25),.clk(clk),.wout(w82_25));
	PE pe82_26(.x(x26),.w(w82_25),.acc(r82_25),.res(r82_26),.clk(clk),.wout(w82_26));
	PE pe82_27(.x(x27),.w(w82_26),.acc(r82_26),.res(r82_27),.clk(clk),.wout(w82_27));
	PE pe82_28(.x(x28),.w(w82_27),.acc(r82_27),.res(r82_28),.clk(clk),.wout(w82_28));
	PE pe82_29(.x(x29),.w(w82_28),.acc(r82_28),.res(r82_29),.clk(clk),.wout(w82_29));
	PE pe82_30(.x(x30),.w(w82_29),.acc(r82_29),.res(r82_30),.clk(clk),.wout(w82_30));
	PE pe82_31(.x(x31),.w(w82_30),.acc(r82_30),.res(r82_31),.clk(clk),.wout(w82_31));
	PE pe82_32(.x(x32),.w(w82_31),.acc(r82_31),.res(r82_32),.clk(clk),.wout(w82_32));
	PE pe82_33(.x(x33),.w(w82_32),.acc(r82_32),.res(r82_33),.clk(clk),.wout(w82_33));
	PE pe82_34(.x(x34),.w(w82_33),.acc(r82_33),.res(r82_34),.clk(clk),.wout(w82_34));
	PE pe82_35(.x(x35),.w(w82_34),.acc(r82_34),.res(r82_35),.clk(clk),.wout(w82_35));
	PE pe82_36(.x(x36),.w(w82_35),.acc(r82_35),.res(r82_36),.clk(clk),.wout(w82_36));
	PE pe82_37(.x(x37),.w(w82_36),.acc(r82_36),.res(r82_37),.clk(clk),.wout(w82_37));
	PE pe82_38(.x(x38),.w(w82_37),.acc(r82_37),.res(r82_38),.clk(clk),.wout(w82_38));
	PE pe82_39(.x(x39),.w(w82_38),.acc(r82_38),.res(r82_39),.clk(clk),.wout(w82_39));
	PE pe82_40(.x(x40),.w(w82_39),.acc(r82_39),.res(r82_40),.clk(clk),.wout(w82_40));
	PE pe82_41(.x(x41),.w(w82_40),.acc(r82_40),.res(r82_41),.clk(clk),.wout(w82_41));
	PE pe82_42(.x(x42),.w(w82_41),.acc(r82_41),.res(r82_42),.clk(clk),.wout(w82_42));
	PE pe82_43(.x(x43),.w(w82_42),.acc(r82_42),.res(r82_43),.clk(clk),.wout(w82_43));
	PE pe82_44(.x(x44),.w(w82_43),.acc(r82_43),.res(r82_44),.clk(clk),.wout(w82_44));
	PE pe82_45(.x(x45),.w(w82_44),.acc(r82_44),.res(r82_45),.clk(clk),.wout(w82_45));
	PE pe82_46(.x(x46),.w(w82_45),.acc(r82_45),.res(r82_46),.clk(clk),.wout(w82_46));
	PE pe82_47(.x(x47),.w(w82_46),.acc(r82_46),.res(r82_47),.clk(clk),.wout(w82_47));
	PE pe82_48(.x(x48),.w(w82_47),.acc(r82_47),.res(r82_48),.clk(clk),.wout(w82_48));
	PE pe82_49(.x(x49),.w(w82_48),.acc(r82_48),.res(r82_49),.clk(clk),.wout(w82_49));
	PE pe82_50(.x(x50),.w(w82_49),.acc(r82_49),.res(r82_50),.clk(clk),.wout(w82_50));
	PE pe82_51(.x(x51),.w(w82_50),.acc(r82_50),.res(r82_51),.clk(clk),.wout(w82_51));
	PE pe82_52(.x(x52),.w(w82_51),.acc(r82_51),.res(r82_52),.clk(clk),.wout(w82_52));
	PE pe82_53(.x(x53),.w(w82_52),.acc(r82_52),.res(r82_53),.clk(clk),.wout(w82_53));
	PE pe82_54(.x(x54),.w(w82_53),.acc(r82_53),.res(r82_54),.clk(clk),.wout(w82_54));
	PE pe82_55(.x(x55),.w(w82_54),.acc(r82_54),.res(r82_55),.clk(clk),.wout(w82_55));
	PE pe82_56(.x(x56),.w(w82_55),.acc(r82_55),.res(r82_56),.clk(clk),.wout(w82_56));
	PE pe82_57(.x(x57),.w(w82_56),.acc(r82_56),.res(r82_57),.clk(clk),.wout(w82_57));
	PE pe82_58(.x(x58),.w(w82_57),.acc(r82_57),.res(r82_58),.clk(clk),.wout(w82_58));
	PE pe82_59(.x(x59),.w(w82_58),.acc(r82_58),.res(r82_59),.clk(clk),.wout(w82_59));
	PE pe82_60(.x(x60),.w(w82_59),.acc(r82_59),.res(r82_60),.clk(clk),.wout(w82_60));
	PE pe82_61(.x(x61),.w(w82_60),.acc(r82_60),.res(r82_61),.clk(clk),.wout(w82_61));
	PE pe82_62(.x(x62),.w(w82_61),.acc(r82_61),.res(r82_62),.clk(clk),.wout(w82_62));
	PE pe82_63(.x(x63),.w(w82_62),.acc(r82_62),.res(r82_63),.clk(clk),.wout(w82_63));
	PE pe82_64(.x(x64),.w(w82_63),.acc(r82_63),.res(r82_64),.clk(clk),.wout(w82_64));
	PE pe82_65(.x(x65),.w(w82_64),.acc(r82_64),.res(r82_65),.clk(clk),.wout(w82_65));
	PE pe82_66(.x(x66),.w(w82_65),.acc(r82_65),.res(r82_66),.clk(clk),.wout(w82_66));
	PE pe82_67(.x(x67),.w(w82_66),.acc(r82_66),.res(r82_67),.clk(clk),.wout(w82_67));
	PE pe82_68(.x(x68),.w(w82_67),.acc(r82_67),.res(r82_68),.clk(clk),.wout(w82_68));
	PE pe82_69(.x(x69),.w(w82_68),.acc(r82_68),.res(r82_69),.clk(clk),.wout(w82_69));
	PE pe82_70(.x(x70),.w(w82_69),.acc(r82_69),.res(r82_70),.clk(clk),.wout(w82_70));
	PE pe82_71(.x(x71),.w(w82_70),.acc(r82_70),.res(r82_71),.clk(clk),.wout(w82_71));
	PE pe82_72(.x(x72),.w(w82_71),.acc(r82_71),.res(r82_72),.clk(clk),.wout(w82_72));
	PE pe82_73(.x(x73),.w(w82_72),.acc(r82_72),.res(r82_73),.clk(clk),.wout(w82_73));
	PE pe82_74(.x(x74),.w(w82_73),.acc(r82_73),.res(r82_74),.clk(clk),.wout(w82_74));
	PE pe82_75(.x(x75),.w(w82_74),.acc(r82_74),.res(r82_75),.clk(clk),.wout(w82_75));
	PE pe82_76(.x(x76),.w(w82_75),.acc(r82_75),.res(r82_76),.clk(clk),.wout(w82_76));
	PE pe82_77(.x(x77),.w(w82_76),.acc(r82_76),.res(r82_77),.clk(clk),.wout(w82_77));
	PE pe82_78(.x(x78),.w(w82_77),.acc(r82_77),.res(r82_78),.clk(clk),.wout(w82_78));
	PE pe82_79(.x(x79),.w(w82_78),.acc(r82_78),.res(r82_79),.clk(clk),.wout(w82_79));
	PE pe82_80(.x(x80),.w(w82_79),.acc(r82_79),.res(r82_80),.clk(clk),.wout(w82_80));
	PE pe82_81(.x(x81),.w(w82_80),.acc(r82_80),.res(r82_81),.clk(clk),.wout(w82_81));
	PE pe82_82(.x(x82),.w(w82_81),.acc(r82_81),.res(r82_82),.clk(clk),.wout(w82_82));
	PE pe82_83(.x(x83),.w(w82_82),.acc(r82_82),.res(r82_83),.clk(clk),.wout(w82_83));
	PE pe82_84(.x(x84),.w(w82_83),.acc(r82_83),.res(r82_84),.clk(clk),.wout(w82_84));
	PE pe82_85(.x(x85),.w(w82_84),.acc(r82_84),.res(r82_85),.clk(clk),.wout(w82_85));
	PE pe82_86(.x(x86),.w(w82_85),.acc(r82_85),.res(r82_86),.clk(clk),.wout(w82_86));
	PE pe82_87(.x(x87),.w(w82_86),.acc(r82_86),.res(r82_87),.clk(clk),.wout(w82_87));
	PE pe82_88(.x(x88),.w(w82_87),.acc(r82_87),.res(r82_88),.clk(clk),.wout(w82_88));
	PE pe82_89(.x(x89),.w(w82_88),.acc(r82_88),.res(r82_89),.clk(clk),.wout(w82_89));
	PE pe82_90(.x(x90),.w(w82_89),.acc(r82_89),.res(r82_90),.clk(clk),.wout(w82_90));
	PE pe82_91(.x(x91),.w(w82_90),.acc(r82_90),.res(r82_91),.clk(clk),.wout(w82_91));
	PE pe82_92(.x(x92),.w(w82_91),.acc(r82_91),.res(r82_92),.clk(clk),.wout(w82_92));
	PE pe82_93(.x(x93),.w(w82_92),.acc(r82_92),.res(r82_93),.clk(clk),.wout(w82_93));
	PE pe82_94(.x(x94),.w(w82_93),.acc(r82_93),.res(r82_94),.clk(clk),.wout(w82_94));
	PE pe82_95(.x(x95),.w(w82_94),.acc(r82_94),.res(r82_95),.clk(clk),.wout(w82_95));
	PE pe82_96(.x(x96),.w(w82_95),.acc(r82_95),.res(r82_96),.clk(clk),.wout(w82_96));
	PE pe82_97(.x(x97),.w(w82_96),.acc(r82_96),.res(r82_97),.clk(clk),.wout(w82_97));
	PE pe82_98(.x(x98),.w(w82_97),.acc(r82_97),.res(r82_98),.clk(clk),.wout(w82_98));
	PE pe82_99(.x(x99),.w(w82_98),.acc(r82_98),.res(r82_99),.clk(clk),.wout(w82_99));
	PE pe82_100(.x(x100),.w(w82_99),.acc(r82_99),.res(r82_100),.clk(clk),.wout(w82_100));
	PE pe82_101(.x(x101),.w(w82_100),.acc(r82_100),.res(r82_101),.clk(clk),.wout(w82_101));
	PE pe82_102(.x(x102),.w(w82_101),.acc(r82_101),.res(r82_102),.clk(clk),.wout(w82_102));
	PE pe82_103(.x(x103),.w(w82_102),.acc(r82_102),.res(r82_103),.clk(clk),.wout(w82_103));
	PE pe82_104(.x(x104),.w(w82_103),.acc(r82_103),.res(r82_104),.clk(clk),.wout(w82_104));
	PE pe82_105(.x(x105),.w(w82_104),.acc(r82_104),.res(r82_105),.clk(clk),.wout(w82_105));
	PE pe82_106(.x(x106),.w(w82_105),.acc(r82_105),.res(r82_106),.clk(clk),.wout(w82_106));
	PE pe82_107(.x(x107),.w(w82_106),.acc(r82_106),.res(r82_107),.clk(clk),.wout(w82_107));
	PE pe82_108(.x(x108),.w(w82_107),.acc(r82_107),.res(r82_108),.clk(clk),.wout(w82_108));
	PE pe82_109(.x(x109),.w(w82_108),.acc(r82_108),.res(r82_109),.clk(clk),.wout(w82_109));
	PE pe82_110(.x(x110),.w(w82_109),.acc(r82_109),.res(r82_110),.clk(clk),.wout(w82_110));
	PE pe82_111(.x(x111),.w(w82_110),.acc(r82_110),.res(r82_111),.clk(clk),.wout(w82_111));
	PE pe82_112(.x(x112),.w(w82_111),.acc(r82_111),.res(r82_112),.clk(clk),.wout(w82_112));
	PE pe82_113(.x(x113),.w(w82_112),.acc(r82_112),.res(r82_113),.clk(clk),.wout(w82_113));
	PE pe82_114(.x(x114),.w(w82_113),.acc(r82_113),.res(r82_114),.clk(clk),.wout(w82_114));
	PE pe82_115(.x(x115),.w(w82_114),.acc(r82_114),.res(r82_115),.clk(clk),.wout(w82_115));
	PE pe82_116(.x(x116),.w(w82_115),.acc(r82_115),.res(r82_116),.clk(clk),.wout(w82_116));
	PE pe82_117(.x(x117),.w(w82_116),.acc(r82_116),.res(r82_117),.clk(clk),.wout(w82_117));
	PE pe82_118(.x(x118),.w(w82_117),.acc(r82_117),.res(r82_118),.clk(clk),.wout(w82_118));
	PE pe82_119(.x(x119),.w(w82_118),.acc(r82_118),.res(r82_119),.clk(clk),.wout(w82_119));
	PE pe82_120(.x(x120),.w(w82_119),.acc(r82_119),.res(r82_120),.clk(clk),.wout(w82_120));
	PE pe82_121(.x(x121),.w(w82_120),.acc(r82_120),.res(r82_121),.clk(clk),.wout(w82_121));
	PE pe82_122(.x(x122),.w(w82_121),.acc(r82_121),.res(r82_122),.clk(clk),.wout(w82_122));
	PE pe82_123(.x(x123),.w(w82_122),.acc(r82_122),.res(r82_123),.clk(clk),.wout(w82_123));
	PE pe82_124(.x(x124),.w(w82_123),.acc(r82_123),.res(r82_124),.clk(clk),.wout(w82_124));
	PE pe82_125(.x(x125),.w(w82_124),.acc(r82_124),.res(r82_125),.clk(clk),.wout(w82_125));
	PE pe82_126(.x(x126),.w(w82_125),.acc(r82_125),.res(r82_126),.clk(clk),.wout(w82_126));
	PE pe82_127(.x(x127),.w(w82_126),.acc(r82_126),.res(result82),.clk(clk),.wout(weight82));

	PE pe83_0(.x(x0),.w(w83),.acc(32'h0),.res(r83_0),.clk(clk),.wout(w83_0));
	PE pe83_1(.x(x1),.w(w83_0),.acc(r83_0),.res(r83_1),.clk(clk),.wout(w83_1));
	PE pe83_2(.x(x2),.w(w83_1),.acc(r83_1),.res(r83_2),.clk(clk),.wout(w83_2));
	PE pe83_3(.x(x3),.w(w83_2),.acc(r83_2),.res(r83_3),.clk(clk),.wout(w83_3));
	PE pe83_4(.x(x4),.w(w83_3),.acc(r83_3),.res(r83_4),.clk(clk),.wout(w83_4));
	PE pe83_5(.x(x5),.w(w83_4),.acc(r83_4),.res(r83_5),.clk(clk),.wout(w83_5));
	PE pe83_6(.x(x6),.w(w83_5),.acc(r83_5),.res(r83_6),.clk(clk),.wout(w83_6));
	PE pe83_7(.x(x7),.w(w83_6),.acc(r83_6),.res(r83_7),.clk(clk),.wout(w83_7));
	PE pe83_8(.x(x8),.w(w83_7),.acc(r83_7),.res(r83_8),.clk(clk),.wout(w83_8));
	PE pe83_9(.x(x9),.w(w83_8),.acc(r83_8),.res(r83_9),.clk(clk),.wout(w83_9));
	PE pe83_10(.x(x10),.w(w83_9),.acc(r83_9),.res(r83_10),.clk(clk),.wout(w83_10));
	PE pe83_11(.x(x11),.w(w83_10),.acc(r83_10),.res(r83_11),.clk(clk),.wout(w83_11));
	PE pe83_12(.x(x12),.w(w83_11),.acc(r83_11),.res(r83_12),.clk(clk),.wout(w83_12));
	PE pe83_13(.x(x13),.w(w83_12),.acc(r83_12),.res(r83_13),.clk(clk),.wout(w83_13));
	PE pe83_14(.x(x14),.w(w83_13),.acc(r83_13),.res(r83_14),.clk(clk),.wout(w83_14));
	PE pe83_15(.x(x15),.w(w83_14),.acc(r83_14),.res(r83_15),.clk(clk),.wout(w83_15));
	PE pe83_16(.x(x16),.w(w83_15),.acc(r83_15),.res(r83_16),.clk(clk),.wout(w83_16));
	PE pe83_17(.x(x17),.w(w83_16),.acc(r83_16),.res(r83_17),.clk(clk),.wout(w83_17));
	PE pe83_18(.x(x18),.w(w83_17),.acc(r83_17),.res(r83_18),.clk(clk),.wout(w83_18));
	PE pe83_19(.x(x19),.w(w83_18),.acc(r83_18),.res(r83_19),.clk(clk),.wout(w83_19));
	PE pe83_20(.x(x20),.w(w83_19),.acc(r83_19),.res(r83_20),.clk(clk),.wout(w83_20));
	PE pe83_21(.x(x21),.w(w83_20),.acc(r83_20),.res(r83_21),.clk(clk),.wout(w83_21));
	PE pe83_22(.x(x22),.w(w83_21),.acc(r83_21),.res(r83_22),.clk(clk),.wout(w83_22));
	PE pe83_23(.x(x23),.w(w83_22),.acc(r83_22),.res(r83_23),.clk(clk),.wout(w83_23));
	PE pe83_24(.x(x24),.w(w83_23),.acc(r83_23),.res(r83_24),.clk(clk),.wout(w83_24));
	PE pe83_25(.x(x25),.w(w83_24),.acc(r83_24),.res(r83_25),.clk(clk),.wout(w83_25));
	PE pe83_26(.x(x26),.w(w83_25),.acc(r83_25),.res(r83_26),.clk(clk),.wout(w83_26));
	PE pe83_27(.x(x27),.w(w83_26),.acc(r83_26),.res(r83_27),.clk(clk),.wout(w83_27));
	PE pe83_28(.x(x28),.w(w83_27),.acc(r83_27),.res(r83_28),.clk(clk),.wout(w83_28));
	PE pe83_29(.x(x29),.w(w83_28),.acc(r83_28),.res(r83_29),.clk(clk),.wout(w83_29));
	PE pe83_30(.x(x30),.w(w83_29),.acc(r83_29),.res(r83_30),.clk(clk),.wout(w83_30));
	PE pe83_31(.x(x31),.w(w83_30),.acc(r83_30),.res(r83_31),.clk(clk),.wout(w83_31));
	PE pe83_32(.x(x32),.w(w83_31),.acc(r83_31),.res(r83_32),.clk(clk),.wout(w83_32));
	PE pe83_33(.x(x33),.w(w83_32),.acc(r83_32),.res(r83_33),.clk(clk),.wout(w83_33));
	PE pe83_34(.x(x34),.w(w83_33),.acc(r83_33),.res(r83_34),.clk(clk),.wout(w83_34));
	PE pe83_35(.x(x35),.w(w83_34),.acc(r83_34),.res(r83_35),.clk(clk),.wout(w83_35));
	PE pe83_36(.x(x36),.w(w83_35),.acc(r83_35),.res(r83_36),.clk(clk),.wout(w83_36));
	PE pe83_37(.x(x37),.w(w83_36),.acc(r83_36),.res(r83_37),.clk(clk),.wout(w83_37));
	PE pe83_38(.x(x38),.w(w83_37),.acc(r83_37),.res(r83_38),.clk(clk),.wout(w83_38));
	PE pe83_39(.x(x39),.w(w83_38),.acc(r83_38),.res(r83_39),.clk(clk),.wout(w83_39));
	PE pe83_40(.x(x40),.w(w83_39),.acc(r83_39),.res(r83_40),.clk(clk),.wout(w83_40));
	PE pe83_41(.x(x41),.w(w83_40),.acc(r83_40),.res(r83_41),.clk(clk),.wout(w83_41));
	PE pe83_42(.x(x42),.w(w83_41),.acc(r83_41),.res(r83_42),.clk(clk),.wout(w83_42));
	PE pe83_43(.x(x43),.w(w83_42),.acc(r83_42),.res(r83_43),.clk(clk),.wout(w83_43));
	PE pe83_44(.x(x44),.w(w83_43),.acc(r83_43),.res(r83_44),.clk(clk),.wout(w83_44));
	PE pe83_45(.x(x45),.w(w83_44),.acc(r83_44),.res(r83_45),.clk(clk),.wout(w83_45));
	PE pe83_46(.x(x46),.w(w83_45),.acc(r83_45),.res(r83_46),.clk(clk),.wout(w83_46));
	PE pe83_47(.x(x47),.w(w83_46),.acc(r83_46),.res(r83_47),.clk(clk),.wout(w83_47));
	PE pe83_48(.x(x48),.w(w83_47),.acc(r83_47),.res(r83_48),.clk(clk),.wout(w83_48));
	PE pe83_49(.x(x49),.w(w83_48),.acc(r83_48),.res(r83_49),.clk(clk),.wout(w83_49));
	PE pe83_50(.x(x50),.w(w83_49),.acc(r83_49),.res(r83_50),.clk(clk),.wout(w83_50));
	PE pe83_51(.x(x51),.w(w83_50),.acc(r83_50),.res(r83_51),.clk(clk),.wout(w83_51));
	PE pe83_52(.x(x52),.w(w83_51),.acc(r83_51),.res(r83_52),.clk(clk),.wout(w83_52));
	PE pe83_53(.x(x53),.w(w83_52),.acc(r83_52),.res(r83_53),.clk(clk),.wout(w83_53));
	PE pe83_54(.x(x54),.w(w83_53),.acc(r83_53),.res(r83_54),.clk(clk),.wout(w83_54));
	PE pe83_55(.x(x55),.w(w83_54),.acc(r83_54),.res(r83_55),.clk(clk),.wout(w83_55));
	PE pe83_56(.x(x56),.w(w83_55),.acc(r83_55),.res(r83_56),.clk(clk),.wout(w83_56));
	PE pe83_57(.x(x57),.w(w83_56),.acc(r83_56),.res(r83_57),.clk(clk),.wout(w83_57));
	PE pe83_58(.x(x58),.w(w83_57),.acc(r83_57),.res(r83_58),.clk(clk),.wout(w83_58));
	PE pe83_59(.x(x59),.w(w83_58),.acc(r83_58),.res(r83_59),.clk(clk),.wout(w83_59));
	PE pe83_60(.x(x60),.w(w83_59),.acc(r83_59),.res(r83_60),.clk(clk),.wout(w83_60));
	PE pe83_61(.x(x61),.w(w83_60),.acc(r83_60),.res(r83_61),.clk(clk),.wout(w83_61));
	PE pe83_62(.x(x62),.w(w83_61),.acc(r83_61),.res(r83_62),.clk(clk),.wout(w83_62));
	PE pe83_63(.x(x63),.w(w83_62),.acc(r83_62),.res(r83_63),.clk(clk),.wout(w83_63));
	PE pe83_64(.x(x64),.w(w83_63),.acc(r83_63),.res(r83_64),.clk(clk),.wout(w83_64));
	PE pe83_65(.x(x65),.w(w83_64),.acc(r83_64),.res(r83_65),.clk(clk),.wout(w83_65));
	PE pe83_66(.x(x66),.w(w83_65),.acc(r83_65),.res(r83_66),.clk(clk),.wout(w83_66));
	PE pe83_67(.x(x67),.w(w83_66),.acc(r83_66),.res(r83_67),.clk(clk),.wout(w83_67));
	PE pe83_68(.x(x68),.w(w83_67),.acc(r83_67),.res(r83_68),.clk(clk),.wout(w83_68));
	PE pe83_69(.x(x69),.w(w83_68),.acc(r83_68),.res(r83_69),.clk(clk),.wout(w83_69));
	PE pe83_70(.x(x70),.w(w83_69),.acc(r83_69),.res(r83_70),.clk(clk),.wout(w83_70));
	PE pe83_71(.x(x71),.w(w83_70),.acc(r83_70),.res(r83_71),.clk(clk),.wout(w83_71));
	PE pe83_72(.x(x72),.w(w83_71),.acc(r83_71),.res(r83_72),.clk(clk),.wout(w83_72));
	PE pe83_73(.x(x73),.w(w83_72),.acc(r83_72),.res(r83_73),.clk(clk),.wout(w83_73));
	PE pe83_74(.x(x74),.w(w83_73),.acc(r83_73),.res(r83_74),.clk(clk),.wout(w83_74));
	PE pe83_75(.x(x75),.w(w83_74),.acc(r83_74),.res(r83_75),.clk(clk),.wout(w83_75));
	PE pe83_76(.x(x76),.w(w83_75),.acc(r83_75),.res(r83_76),.clk(clk),.wout(w83_76));
	PE pe83_77(.x(x77),.w(w83_76),.acc(r83_76),.res(r83_77),.clk(clk),.wout(w83_77));
	PE pe83_78(.x(x78),.w(w83_77),.acc(r83_77),.res(r83_78),.clk(clk),.wout(w83_78));
	PE pe83_79(.x(x79),.w(w83_78),.acc(r83_78),.res(r83_79),.clk(clk),.wout(w83_79));
	PE pe83_80(.x(x80),.w(w83_79),.acc(r83_79),.res(r83_80),.clk(clk),.wout(w83_80));
	PE pe83_81(.x(x81),.w(w83_80),.acc(r83_80),.res(r83_81),.clk(clk),.wout(w83_81));
	PE pe83_82(.x(x82),.w(w83_81),.acc(r83_81),.res(r83_82),.clk(clk),.wout(w83_82));
	PE pe83_83(.x(x83),.w(w83_82),.acc(r83_82),.res(r83_83),.clk(clk),.wout(w83_83));
	PE pe83_84(.x(x84),.w(w83_83),.acc(r83_83),.res(r83_84),.clk(clk),.wout(w83_84));
	PE pe83_85(.x(x85),.w(w83_84),.acc(r83_84),.res(r83_85),.clk(clk),.wout(w83_85));
	PE pe83_86(.x(x86),.w(w83_85),.acc(r83_85),.res(r83_86),.clk(clk),.wout(w83_86));
	PE pe83_87(.x(x87),.w(w83_86),.acc(r83_86),.res(r83_87),.clk(clk),.wout(w83_87));
	PE pe83_88(.x(x88),.w(w83_87),.acc(r83_87),.res(r83_88),.clk(clk),.wout(w83_88));
	PE pe83_89(.x(x89),.w(w83_88),.acc(r83_88),.res(r83_89),.clk(clk),.wout(w83_89));
	PE pe83_90(.x(x90),.w(w83_89),.acc(r83_89),.res(r83_90),.clk(clk),.wout(w83_90));
	PE pe83_91(.x(x91),.w(w83_90),.acc(r83_90),.res(r83_91),.clk(clk),.wout(w83_91));
	PE pe83_92(.x(x92),.w(w83_91),.acc(r83_91),.res(r83_92),.clk(clk),.wout(w83_92));
	PE pe83_93(.x(x93),.w(w83_92),.acc(r83_92),.res(r83_93),.clk(clk),.wout(w83_93));
	PE pe83_94(.x(x94),.w(w83_93),.acc(r83_93),.res(r83_94),.clk(clk),.wout(w83_94));
	PE pe83_95(.x(x95),.w(w83_94),.acc(r83_94),.res(r83_95),.clk(clk),.wout(w83_95));
	PE pe83_96(.x(x96),.w(w83_95),.acc(r83_95),.res(r83_96),.clk(clk),.wout(w83_96));
	PE pe83_97(.x(x97),.w(w83_96),.acc(r83_96),.res(r83_97),.clk(clk),.wout(w83_97));
	PE pe83_98(.x(x98),.w(w83_97),.acc(r83_97),.res(r83_98),.clk(clk),.wout(w83_98));
	PE pe83_99(.x(x99),.w(w83_98),.acc(r83_98),.res(r83_99),.clk(clk),.wout(w83_99));
	PE pe83_100(.x(x100),.w(w83_99),.acc(r83_99),.res(r83_100),.clk(clk),.wout(w83_100));
	PE pe83_101(.x(x101),.w(w83_100),.acc(r83_100),.res(r83_101),.clk(clk),.wout(w83_101));
	PE pe83_102(.x(x102),.w(w83_101),.acc(r83_101),.res(r83_102),.clk(clk),.wout(w83_102));
	PE pe83_103(.x(x103),.w(w83_102),.acc(r83_102),.res(r83_103),.clk(clk),.wout(w83_103));
	PE pe83_104(.x(x104),.w(w83_103),.acc(r83_103),.res(r83_104),.clk(clk),.wout(w83_104));
	PE pe83_105(.x(x105),.w(w83_104),.acc(r83_104),.res(r83_105),.clk(clk),.wout(w83_105));
	PE pe83_106(.x(x106),.w(w83_105),.acc(r83_105),.res(r83_106),.clk(clk),.wout(w83_106));
	PE pe83_107(.x(x107),.w(w83_106),.acc(r83_106),.res(r83_107),.clk(clk),.wout(w83_107));
	PE pe83_108(.x(x108),.w(w83_107),.acc(r83_107),.res(r83_108),.clk(clk),.wout(w83_108));
	PE pe83_109(.x(x109),.w(w83_108),.acc(r83_108),.res(r83_109),.clk(clk),.wout(w83_109));
	PE pe83_110(.x(x110),.w(w83_109),.acc(r83_109),.res(r83_110),.clk(clk),.wout(w83_110));
	PE pe83_111(.x(x111),.w(w83_110),.acc(r83_110),.res(r83_111),.clk(clk),.wout(w83_111));
	PE pe83_112(.x(x112),.w(w83_111),.acc(r83_111),.res(r83_112),.clk(clk),.wout(w83_112));
	PE pe83_113(.x(x113),.w(w83_112),.acc(r83_112),.res(r83_113),.clk(clk),.wout(w83_113));
	PE pe83_114(.x(x114),.w(w83_113),.acc(r83_113),.res(r83_114),.clk(clk),.wout(w83_114));
	PE pe83_115(.x(x115),.w(w83_114),.acc(r83_114),.res(r83_115),.clk(clk),.wout(w83_115));
	PE pe83_116(.x(x116),.w(w83_115),.acc(r83_115),.res(r83_116),.clk(clk),.wout(w83_116));
	PE pe83_117(.x(x117),.w(w83_116),.acc(r83_116),.res(r83_117),.clk(clk),.wout(w83_117));
	PE pe83_118(.x(x118),.w(w83_117),.acc(r83_117),.res(r83_118),.clk(clk),.wout(w83_118));
	PE pe83_119(.x(x119),.w(w83_118),.acc(r83_118),.res(r83_119),.clk(clk),.wout(w83_119));
	PE pe83_120(.x(x120),.w(w83_119),.acc(r83_119),.res(r83_120),.clk(clk),.wout(w83_120));
	PE pe83_121(.x(x121),.w(w83_120),.acc(r83_120),.res(r83_121),.clk(clk),.wout(w83_121));
	PE pe83_122(.x(x122),.w(w83_121),.acc(r83_121),.res(r83_122),.clk(clk),.wout(w83_122));
	PE pe83_123(.x(x123),.w(w83_122),.acc(r83_122),.res(r83_123),.clk(clk),.wout(w83_123));
	PE pe83_124(.x(x124),.w(w83_123),.acc(r83_123),.res(r83_124),.clk(clk),.wout(w83_124));
	PE pe83_125(.x(x125),.w(w83_124),.acc(r83_124),.res(r83_125),.clk(clk),.wout(w83_125));
	PE pe83_126(.x(x126),.w(w83_125),.acc(r83_125),.res(r83_126),.clk(clk),.wout(w83_126));
	PE pe83_127(.x(x127),.w(w83_126),.acc(r83_126),.res(result83),.clk(clk),.wout(weight83));

	PE pe84_0(.x(x0),.w(w84),.acc(32'h0),.res(r84_0),.clk(clk),.wout(w84_0));
	PE pe84_1(.x(x1),.w(w84_0),.acc(r84_0),.res(r84_1),.clk(clk),.wout(w84_1));
	PE pe84_2(.x(x2),.w(w84_1),.acc(r84_1),.res(r84_2),.clk(clk),.wout(w84_2));
	PE pe84_3(.x(x3),.w(w84_2),.acc(r84_2),.res(r84_3),.clk(clk),.wout(w84_3));
	PE pe84_4(.x(x4),.w(w84_3),.acc(r84_3),.res(r84_4),.clk(clk),.wout(w84_4));
	PE pe84_5(.x(x5),.w(w84_4),.acc(r84_4),.res(r84_5),.clk(clk),.wout(w84_5));
	PE pe84_6(.x(x6),.w(w84_5),.acc(r84_5),.res(r84_6),.clk(clk),.wout(w84_6));
	PE pe84_7(.x(x7),.w(w84_6),.acc(r84_6),.res(r84_7),.clk(clk),.wout(w84_7));
	PE pe84_8(.x(x8),.w(w84_7),.acc(r84_7),.res(r84_8),.clk(clk),.wout(w84_8));
	PE pe84_9(.x(x9),.w(w84_8),.acc(r84_8),.res(r84_9),.clk(clk),.wout(w84_9));
	PE pe84_10(.x(x10),.w(w84_9),.acc(r84_9),.res(r84_10),.clk(clk),.wout(w84_10));
	PE pe84_11(.x(x11),.w(w84_10),.acc(r84_10),.res(r84_11),.clk(clk),.wout(w84_11));
	PE pe84_12(.x(x12),.w(w84_11),.acc(r84_11),.res(r84_12),.clk(clk),.wout(w84_12));
	PE pe84_13(.x(x13),.w(w84_12),.acc(r84_12),.res(r84_13),.clk(clk),.wout(w84_13));
	PE pe84_14(.x(x14),.w(w84_13),.acc(r84_13),.res(r84_14),.clk(clk),.wout(w84_14));
	PE pe84_15(.x(x15),.w(w84_14),.acc(r84_14),.res(r84_15),.clk(clk),.wout(w84_15));
	PE pe84_16(.x(x16),.w(w84_15),.acc(r84_15),.res(r84_16),.clk(clk),.wout(w84_16));
	PE pe84_17(.x(x17),.w(w84_16),.acc(r84_16),.res(r84_17),.clk(clk),.wout(w84_17));
	PE pe84_18(.x(x18),.w(w84_17),.acc(r84_17),.res(r84_18),.clk(clk),.wout(w84_18));
	PE pe84_19(.x(x19),.w(w84_18),.acc(r84_18),.res(r84_19),.clk(clk),.wout(w84_19));
	PE pe84_20(.x(x20),.w(w84_19),.acc(r84_19),.res(r84_20),.clk(clk),.wout(w84_20));
	PE pe84_21(.x(x21),.w(w84_20),.acc(r84_20),.res(r84_21),.clk(clk),.wout(w84_21));
	PE pe84_22(.x(x22),.w(w84_21),.acc(r84_21),.res(r84_22),.clk(clk),.wout(w84_22));
	PE pe84_23(.x(x23),.w(w84_22),.acc(r84_22),.res(r84_23),.clk(clk),.wout(w84_23));
	PE pe84_24(.x(x24),.w(w84_23),.acc(r84_23),.res(r84_24),.clk(clk),.wout(w84_24));
	PE pe84_25(.x(x25),.w(w84_24),.acc(r84_24),.res(r84_25),.clk(clk),.wout(w84_25));
	PE pe84_26(.x(x26),.w(w84_25),.acc(r84_25),.res(r84_26),.clk(clk),.wout(w84_26));
	PE pe84_27(.x(x27),.w(w84_26),.acc(r84_26),.res(r84_27),.clk(clk),.wout(w84_27));
	PE pe84_28(.x(x28),.w(w84_27),.acc(r84_27),.res(r84_28),.clk(clk),.wout(w84_28));
	PE pe84_29(.x(x29),.w(w84_28),.acc(r84_28),.res(r84_29),.clk(clk),.wout(w84_29));
	PE pe84_30(.x(x30),.w(w84_29),.acc(r84_29),.res(r84_30),.clk(clk),.wout(w84_30));
	PE pe84_31(.x(x31),.w(w84_30),.acc(r84_30),.res(r84_31),.clk(clk),.wout(w84_31));
	PE pe84_32(.x(x32),.w(w84_31),.acc(r84_31),.res(r84_32),.clk(clk),.wout(w84_32));
	PE pe84_33(.x(x33),.w(w84_32),.acc(r84_32),.res(r84_33),.clk(clk),.wout(w84_33));
	PE pe84_34(.x(x34),.w(w84_33),.acc(r84_33),.res(r84_34),.clk(clk),.wout(w84_34));
	PE pe84_35(.x(x35),.w(w84_34),.acc(r84_34),.res(r84_35),.clk(clk),.wout(w84_35));
	PE pe84_36(.x(x36),.w(w84_35),.acc(r84_35),.res(r84_36),.clk(clk),.wout(w84_36));
	PE pe84_37(.x(x37),.w(w84_36),.acc(r84_36),.res(r84_37),.clk(clk),.wout(w84_37));
	PE pe84_38(.x(x38),.w(w84_37),.acc(r84_37),.res(r84_38),.clk(clk),.wout(w84_38));
	PE pe84_39(.x(x39),.w(w84_38),.acc(r84_38),.res(r84_39),.clk(clk),.wout(w84_39));
	PE pe84_40(.x(x40),.w(w84_39),.acc(r84_39),.res(r84_40),.clk(clk),.wout(w84_40));
	PE pe84_41(.x(x41),.w(w84_40),.acc(r84_40),.res(r84_41),.clk(clk),.wout(w84_41));
	PE pe84_42(.x(x42),.w(w84_41),.acc(r84_41),.res(r84_42),.clk(clk),.wout(w84_42));
	PE pe84_43(.x(x43),.w(w84_42),.acc(r84_42),.res(r84_43),.clk(clk),.wout(w84_43));
	PE pe84_44(.x(x44),.w(w84_43),.acc(r84_43),.res(r84_44),.clk(clk),.wout(w84_44));
	PE pe84_45(.x(x45),.w(w84_44),.acc(r84_44),.res(r84_45),.clk(clk),.wout(w84_45));
	PE pe84_46(.x(x46),.w(w84_45),.acc(r84_45),.res(r84_46),.clk(clk),.wout(w84_46));
	PE pe84_47(.x(x47),.w(w84_46),.acc(r84_46),.res(r84_47),.clk(clk),.wout(w84_47));
	PE pe84_48(.x(x48),.w(w84_47),.acc(r84_47),.res(r84_48),.clk(clk),.wout(w84_48));
	PE pe84_49(.x(x49),.w(w84_48),.acc(r84_48),.res(r84_49),.clk(clk),.wout(w84_49));
	PE pe84_50(.x(x50),.w(w84_49),.acc(r84_49),.res(r84_50),.clk(clk),.wout(w84_50));
	PE pe84_51(.x(x51),.w(w84_50),.acc(r84_50),.res(r84_51),.clk(clk),.wout(w84_51));
	PE pe84_52(.x(x52),.w(w84_51),.acc(r84_51),.res(r84_52),.clk(clk),.wout(w84_52));
	PE pe84_53(.x(x53),.w(w84_52),.acc(r84_52),.res(r84_53),.clk(clk),.wout(w84_53));
	PE pe84_54(.x(x54),.w(w84_53),.acc(r84_53),.res(r84_54),.clk(clk),.wout(w84_54));
	PE pe84_55(.x(x55),.w(w84_54),.acc(r84_54),.res(r84_55),.clk(clk),.wout(w84_55));
	PE pe84_56(.x(x56),.w(w84_55),.acc(r84_55),.res(r84_56),.clk(clk),.wout(w84_56));
	PE pe84_57(.x(x57),.w(w84_56),.acc(r84_56),.res(r84_57),.clk(clk),.wout(w84_57));
	PE pe84_58(.x(x58),.w(w84_57),.acc(r84_57),.res(r84_58),.clk(clk),.wout(w84_58));
	PE pe84_59(.x(x59),.w(w84_58),.acc(r84_58),.res(r84_59),.clk(clk),.wout(w84_59));
	PE pe84_60(.x(x60),.w(w84_59),.acc(r84_59),.res(r84_60),.clk(clk),.wout(w84_60));
	PE pe84_61(.x(x61),.w(w84_60),.acc(r84_60),.res(r84_61),.clk(clk),.wout(w84_61));
	PE pe84_62(.x(x62),.w(w84_61),.acc(r84_61),.res(r84_62),.clk(clk),.wout(w84_62));
	PE pe84_63(.x(x63),.w(w84_62),.acc(r84_62),.res(r84_63),.clk(clk),.wout(w84_63));
	PE pe84_64(.x(x64),.w(w84_63),.acc(r84_63),.res(r84_64),.clk(clk),.wout(w84_64));
	PE pe84_65(.x(x65),.w(w84_64),.acc(r84_64),.res(r84_65),.clk(clk),.wout(w84_65));
	PE pe84_66(.x(x66),.w(w84_65),.acc(r84_65),.res(r84_66),.clk(clk),.wout(w84_66));
	PE pe84_67(.x(x67),.w(w84_66),.acc(r84_66),.res(r84_67),.clk(clk),.wout(w84_67));
	PE pe84_68(.x(x68),.w(w84_67),.acc(r84_67),.res(r84_68),.clk(clk),.wout(w84_68));
	PE pe84_69(.x(x69),.w(w84_68),.acc(r84_68),.res(r84_69),.clk(clk),.wout(w84_69));
	PE pe84_70(.x(x70),.w(w84_69),.acc(r84_69),.res(r84_70),.clk(clk),.wout(w84_70));
	PE pe84_71(.x(x71),.w(w84_70),.acc(r84_70),.res(r84_71),.clk(clk),.wout(w84_71));
	PE pe84_72(.x(x72),.w(w84_71),.acc(r84_71),.res(r84_72),.clk(clk),.wout(w84_72));
	PE pe84_73(.x(x73),.w(w84_72),.acc(r84_72),.res(r84_73),.clk(clk),.wout(w84_73));
	PE pe84_74(.x(x74),.w(w84_73),.acc(r84_73),.res(r84_74),.clk(clk),.wout(w84_74));
	PE pe84_75(.x(x75),.w(w84_74),.acc(r84_74),.res(r84_75),.clk(clk),.wout(w84_75));
	PE pe84_76(.x(x76),.w(w84_75),.acc(r84_75),.res(r84_76),.clk(clk),.wout(w84_76));
	PE pe84_77(.x(x77),.w(w84_76),.acc(r84_76),.res(r84_77),.clk(clk),.wout(w84_77));
	PE pe84_78(.x(x78),.w(w84_77),.acc(r84_77),.res(r84_78),.clk(clk),.wout(w84_78));
	PE pe84_79(.x(x79),.w(w84_78),.acc(r84_78),.res(r84_79),.clk(clk),.wout(w84_79));
	PE pe84_80(.x(x80),.w(w84_79),.acc(r84_79),.res(r84_80),.clk(clk),.wout(w84_80));
	PE pe84_81(.x(x81),.w(w84_80),.acc(r84_80),.res(r84_81),.clk(clk),.wout(w84_81));
	PE pe84_82(.x(x82),.w(w84_81),.acc(r84_81),.res(r84_82),.clk(clk),.wout(w84_82));
	PE pe84_83(.x(x83),.w(w84_82),.acc(r84_82),.res(r84_83),.clk(clk),.wout(w84_83));
	PE pe84_84(.x(x84),.w(w84_83),.acc(r84_83),.res(r84_84),.clk(clk),.wout(w84_84));
	PE pe84_85(.x(x85),.w(w84_84),.acc(r84_84),.res(r84_85),.clk(clk),.wout(w84_85));
	PE pe84_86(.x(x86),.w(w84_85),.acc(r84_85),.res(r84_86),.clk(clk),.wout(w84_86));
	PE pe84_87(.x(x87),.w(w84_86),.acc(r84_86),.res(r84_87),.clk(clk),.wout(w84_87));
	PE pe84_88(.x(x88),.w(w84_87),.acc(r84_87),.res(r84_88),.clk(clk),.wout(w84_88));
	PE pe84_89(.x(x89),.w(w84_88),.acc(r84_88),.res(r84_89),.clk(clk),.wout(w84_89));
	PE pe84_90(.x(x90),.w(w84_89),.acc(r84_89),.res(r84_90),.clk(clk),.wout(w84_90));
	PE pe84_91(.x(x91),.w(w84_90),.acc(r84_90),.res(r84_91),.clk(clk),.wout(w84_91));
	PE pe84_92(.x(x92),.w(w84_91),.acc(r84_91),.res(r84_92),.clk(clk),.wout(w84_92));
	PE pe84_93(.x(x93),.w(w84_92),.acc(r84_92),.res(r84_93),.clk(clk),.wout(w84_93));
	PE pe84_94(.x(x94),.w(w84_93),.acc(r84_93),.res(r84_94),.clk(clk),.wout(w84_94));
	PE pe84_95(.x(x95),.w(w84_94),.acc(r84_94),.res(r84_95),.clk(clk),.wout(w84_95));
	PE pe84_96(.x(x96),.w(w84_95),.acc(r84_95),.res(r84_96),.clk(clk),.wout(w84_96));
	PE pe84_97(.x(x97),.w(w84_96),.acc(r84_96),.res(r84_97),.clk(clk),.wout(w84_97));
	PE pe84_98(.x(x98),.w(w84_97),.acc(r84_97),.res(r84_98),.clk(clk),.wout(w84_98));
	PE pe84_99(.x(x99),.w(w84_98),.acc(r84_98),.res(r84_99),.clk(clk),.wout(w84_99));
	PE pe84_100(.x(x100),.w(w84_99),.acc(r84_99),.res(r84_100),.clk(clk),.wout(w84_100));
	PE pe84_101(.x(x101),.w(w84_100),.acc(r84_100),.res(r84_101),.clk(clk),.wout(w84_101));
	PE pe84_102(.x(x102),.w(w84_101),.acc(r84_101),.res(r84_102),.clk(clk),.wout(w84_102));
	PE pe84_103(.x(x103),.w(w84_102),.acc(r84_102),.res(r84_103),.clk(clk),.wout(w84_103));
	PE pe84_104(.x(x104),.w(w84_103),.acc(r84_103),.res(r84_104),.clk(clk),.wout(w84_104));
	PE pe84_105(.x(x105),.w(w84_104),.acc(r84_104),.res(r84_105),.clk(clk),.wout(w84_105));
	PE pe84_106(.x(x106),.w(w84_105),.acc(r84_105),.res(r84_106),.clk(clk),.wout(w84_106));
	PE pe84_107(.x(x107),.w(w84_106),.acc(r84_106),.res(r84_107),.clk(clk),.wout(w84_107));
	PE pe84_108(.x(x108),.w(w84_107),.acc(r84_107),.res(r84_108),.clk(clk),.wout(w84_108));
	PE pe84_109(.x(x109),.w(w84_108),.acc(r84_108),.res(r84_109),.clk(clk),.wout(w84_109));
	PE pe84_110(.x(x110),.w(w84_109),.acc(r84_109),.res(r84_110),.clk(clk),.wout(w84_110));
	PE pe84_111(.x(x111),.w(w84_110),.acc(r84_110),.res(r84_111),.clk(clk),.wout(w84_111));
	PE pe84_112(.x(x112),.w(w84_111),.acc(r84_111),.res(r84_112),.clk(clk),.wout(w84_112));
	PE pe84_113(.x(x113),.w(w84_112),.acc(r84_112),.res(r84_113),.clk(clk),.wout(w84_113));
	PE pe84_114(.x(x114),.w(w84_113),.acc(r84_113),.res(r84_114),.clk(clk),.wout(w84_114));
	PE pe84_115(.x(x115),.w(w84_114),.acc(r84_114),.res(r84_115),.clk(clk),.wout(w84_115));
	PE pe84_116(.x(x116),.w(w84_115),.acc(r84_115),.res(r84_116),.clk(clk),.wout(w84_116));
	PE pe84_117(.x(x117),.w(w84_116),.acc(r84_116),.res(r84_117),.clk(clk),.wout(w84_117));
	PE pe84_118(.x(x118),.w(w84_117),.acc(r84_117),.res(r84_118),.clk(clk),.wout(w84_118));
	PE pe84_119(.x(x119),.w(w84_118),.acc(r84_118),.res(r84_119),.clk(clk),.wout(w84_119));
	PE pe84_120(.x(x120),.w(w84_119),.acc(r84_119),.res(r84_120),.clk(clk),.wout(w84_120));
	PE pe84_121(.x(x121),.w(w84_120),.acc(r84_120),.res(r84_121),.clk(clk),.wout(w84_121));
	PE pe84_122(.x(x122),.w(w84_121),.acc(r84_121),.res(r84_122),.clk(clk),.wout(w84_122));
	PE pe84_123(.x(x123),.w(w84_122),.acc(r84_122),.res(r84_123),.clk(clk),.wout(w84_123));
	PE pe84_124(.x(x124),.w(w84_123),.acc(r84_123),.res(r84_124),.clk(clk),.wout(w84_124));
	PE pe84_125(.x(x125),.w(w84_124),.acc(r84_124),.res(r84_125),.clk(clk),.wout(w84_125));
	PE pe84_126(.x(x126),.w(w84_125),.acc(r84_125),.res(r84_126),.clk(clk),.wout(w84_126));
	PE pe84_127(.x(x127),.w(w84_126),.acc(r84_126),.res(result84),.clk(clk),.wout(weight84));

	PE pe85_0(.x(x0),.w(w85),.acc(32'h0),.res(r85_0),.clk(clk),.wout(w85_0));
	PE pe85_1(.x(x1),.w(w85_0),.acc(r85_0),.res(r85_1),.clk(clk),.wout(w85_1));
	PE pe85_2(.x(x2),.w(w85_1),.acc(r85_1),.res(r85_2),.clk(clk),.wout(w85_2));
	PE pe85_3(.x(x3),.w(w85_2),.acc(r85_2),.res(r85_3),.clk(clk),.wout(w85_3));
	PE pe85_4(.x(x4),.w(w85_3),.acc(r85_3),.res(r85_4),.clk(clk),.wout(w85_4));
	PE pe85_5(.x(x5),.w(w85_4),.acc(r85_4),.res(r85_5),.clk(clk),.wout(w85_5));
	PE pe85_6(.x(x6),.w(w85_5),.acc(r85_5),.res(r85_6),.clk(clk),.wout(w85_6));
	PE pe85_7(.x(x7),.w(w85_6),.acc(r85_6),.res(r85_7),.clk(clk),.wout(w85_7));
	PE pe85_8(.x(x8),.w(w85_7),.acc(r85_7),.res(r85_8),.clk(clk),.wout(w85_8));
	PE pe85_9(.x(x9),.w(w85_8),.acc(r85_8),.res(r85_9),.clk(clk),.wout(w85_9));
	PE pe85_10(.x(x10),.w(w85_9),.acc(r85_9),.res(r85_10),.clk(clk),.wout(w85_10));
	PE pe85_11(.x(x11),.w(w85_10),.acc(r85_10),.res(r85_11),.clk(clk),.wout(w85_11));
	PE pe85_12(.x(x12),.w(w85_11),.acc(r85_11),.res(r85_12),.clk(clk),.wout(w85_12));
	PE pe85_13(.x(x13),.w(w85_12),.acc(r85_12),.res(r85_13),.clk(clk),.wout(w85_13));
	PE pe85_14(.x(x14),.w(w85_13),.acc(r85_13),.res(r85_14),.clk(clk),.wout(w85_14));
	PE pe85_15(.x(x15),.w(w85_14),.acc(r85_14),.res(r85_15),.clk(clk),.wout(w85_15));
	PE pe85_16(.x(x16),.w(w85_15),.acc(r85_15),.res(r85_16),.clk(clk),.wout(w85_16));
	PE pe85_17(.x(x17),.w(w85_16),.acc(r85_16),.res(r85_17),.clk(clk),.wout(w85_17));
	PE pe85_18(.x(x18),.w(w85_17),.acc(r85_17),.res(r85_18),.clk(clk),.wout(w85_18));
	PE pe85_19(.x(x19),.w(w85_18),.acc(r85_18),.res(r85_19),.clk(clk),.wout(w85_19));
	PE pe85_20(.x(x20),.w(w85_19),.acc(r85_19),.res(r85_20),.clk(clk),.wout(w85_20));
	PE pe85_21(.x(x21),.w(w85_20),.acc(r85_20),.res(r85_21),.clk(clk),.wout(w85_21));
	PE pe85_22(.x(x22),.w(w85_21),.acc(r85_21),.res(r85_22),.clk(clk),.wout(w85_22));
	PE pe85_23(.x(x23),.w(w85_22),.acc(r85_22),.res(r85_23),.clk(clk),.wout(w85_23));
	PE pe85_24(.x(x24),.w(w85_23),.acc(r85_23),.res(r85_24),.clk(clk),.wout(w85_24));
	PE pe85_25(.x(x25),.w(w85_24),.acc(r85_24),.res(r85_25),.clk(clk),.wout(w85_25));
	PE pe85_26(.x(x26),.w(w85_25),.acc(r85_25),.res(r85_26),.clk(clk),.wout(w85_26));
	PE pe85_27(.x(x27),.w(w85_26),.acc(r85_26),.res(r85_27),.clk(clk),.wout(w85_27));
	PE pe85_28(.x(x28),.w(w85_27),.acc(r85_27),.res(r85_28),.clk(clk),.wout(w85_28));
	PE pe85_29(.x(x29),.w(w85_28),.acc(r85_28),.res(r85_29),.clk(clk),.wout(w85_29));
	PE pe85_30(.x(x30),.w(w85_29),.acc(r85_29),.res(r85_30),.clk(clk),.wout(w85_30));
	PE pe85_31(.x(x31),.w(w85_30),.acc(r85_30),.res(r85_31),.clk(clk),.wout(w85_31));
	PE pe85_32(.x(x32),.w(w85_31),.acc(r85_31),.res(r85_32),.clk(clk),.wout(w85_32));
	PE pe85_33(.x(x33),.w(w85_32),.acc(r85_32),.res(r85_33),.clk(clk),.wout(w85_33));
	PE pe85_34(.x(x34),.w(w85_33),.acc(r85_33),.res(r85_34),.clk(clk),.wout(w85_34));
	PE pe85_35(.x(x35),.w(w85_34),.acc(r85_34),.res(r85_35),.clk(clk),.wout(w85_35));
	PE pe85_36(.x(x36),.w(w85_35),.acc(r85_35),.res(r85_36),.clk(clk),.wout(w85_36));
	PE pe85_37(.x(x37),.w(w85_36),.acc(r85_36),.res(r85_37),.clk(clk),.wout(w85_37));
	PE pe85_38(.x(x38),.w(w85_37),.acc(r85_37),.res(r85_38),.clk(clk),.wout(w85_38));
	PE pe85_39(.x(x39),.w(w85_38),.acc(r85_38),.res(r85_39),.clk(clk),.wout(w85_39));
	PE pe85_40(.x(x40),.w(w85_39),.acc(r85_39),.res(r85_40),.clk(clk),.wout(w85_40));
	PE pe85_41(.x(x41),.w(w85_40),.acc(r85_40),.res(r85_41),.clk(clk),.wout(w85_41));
	PE pe85_42(.x(x42),.w(w85_41),.acc(r85_41),.res(r85_42),.clk(clk),.wout(w85_42));
	PE pe85_43(.x(x43),.w(w85_42),.acc(r85_42),.res(r85_43),.clk(clk),.wout(w85_43));
	PE pe85_44(.x(x44),.w(w85_43),.acc(r85_43),.res(r85_44),.clk(clk),.wout(w85_44));
	PE pe85_45(.x(x45),.w(w85_44),.acc(r85_44),.res(r85_45),.clk(clk),.wout(w85_45));
	PE pe85_46(.x(x46),.w(w85_45),.acc(r85_45),.res(r85_46),.clk(clk),.wout(w85_46));
	PE pe85_47(.x(x47),.w(w85_46),.acc(r85_46),.res(r85_47),.clk(clk),.wout(w85_47));
	PE pe85_48(.x(x48),.w(w85_47),.acc(r85_47),.res(r85_48),.clk(clk),.wout(w85_48));
	PE pe85_49(.x(x49),.w(w85_48),.acc(r85_48),.res(r85_49),.clk(clk),.wout(w85_49));
	PE pe85_50(.x(x50),.w(w85_49),.acc(r85_49),.res(r85_50),.clk(clk),.wout(w85_50));
	PE pe85_51(.x(x51),.w(w85_50),.acc(r85_50),.res(r85_51),.clk(clk),.wout(w85_51));
	PE pe85_52(.x(x52),.w(w85_51),.acc(r85_51),.res(r85_52),.clk(clk),.wout(w85_52));
	PE pe85_53(.x(x53),.w(w85_52),.acc(r85_52),.res(r85_53),.clk(clk),.wout(w85_53));
	PE pe85_54(.x(x54),.w(w85_53),.acc(r85_53),.res(r85_54),.clk(clk),.wout(w85_54));
	PE pe85_55(.x(x55),.w(w85_54),.acc(r85_54),.res(r85_55),.clk(clk),.wout(w85_55));
	PE pe85_56(.x(x56),.w(w85_55),.acc(r85_55),.res(r85_56),.clk(clk),.wout(w85_56));
	PE pe85_57(.x(x57),.w(w85_56),.acc(r85_56),.res(r85_57),.clk(clk),.wout(w85_57));
	PE pe85_58(.x(x58),.w(w85_57),.acc(r85_57),.res(r85_58),.clk(clk),.wout(w85_58));
	PE pe85_59(.x(x59),.w(w85_58),.acc(r85_58),.res(r85_59),.clk(clk),.wout(w85_59));
	PE pe85_60(.x(x60),.w(w85_59),.acc(r85_59),.res(r85_60),.clk(clk),.wout(w85_60));
	PE pe85_61(.x(x61),.w(w85_60),.acc(r85_60),.res(r85_61),.clk(clk),.wout(w85_61));
	PE pe85_62(.x(x62),.w(w85_61),.acc(r85_61),.res(r85_62),.clk(clk),.wout(w85_62));
	PE pe85_63(.x(x63),.w(w85_62),.acc(r85_62),.res(r85_63),.clk(clk),.wout(w85_63));
	PE pe85_64(.x(x64),.w(w85_63),.acc(r85_63),.res(r85_64),.clk(clk),.wout(w85_64));
	PE pe85_65(.x(x65),.w(w85_64),.acc(r85_64),.res(r85_65),.clk(clk),.wout(w85_65));
	PE pe85_66(.x(x66),.w(w85_65),.acc(r85_65),.res(r85_66),.clk(clk),.wout(w85_66));
	PE pe85_67(.x(x67),.w(w85_66),.acc(r85_66),.res(r85_67),.clk(clk),.wout(w85_67));
	PE pe85_68(.x(x68),.w(w85_67),.acc(r85_67),.res(r85_68),.clk(clk),.wout(w85_68));
	PE pe85_69(.x(x69),.w(w85_68),.acc(r85_68),.res(r85_69),.clk(clk),.wout(w85_69));
	PE pe85_70(.x(x70),.w(w85_69),.acc(r85_69),.res(r85_70),.clk(clk),.wout(w85_70));
	PE pe85_71(.x(x71),.w(w85_70),.acc(r85_70),.res(r85_71),.clk(clk),.wout(w85_71));
	PE pe85_72(.x(x72),.w(w85_71),.acc(r85_71),.res(r85_72),.clk(clk),.wout(w85_72));
	PE pe85_73(.x(x73),.w(w85_72),.acc(r85_72),.res(r85_73),.clk(clk),.wout(w85_73));
	PE pe85_74(.x(x74),.w(w85_73),.acc(r85_73),.res(r85_74),.clk(clk),.wout(w85_74));
	PE pe85_75(.x(x75),.w(w85_74),.acc(r85_74),.res(r85_75),.clk(clk),.wout(w85_75));
	PE pe85_76(.x(x76),.w(w85_75),.acc(r85_75),.res(r85_76),.clk(clk),.wout(w85_76));
	PE pe85_77(.x(x77),.w(w85_76),.acc(r85_76),.res(r85_77),.clk(clk),.wout(w85_77));
	PE pe85_78(.x(x78),.w(w85_77),.acc(r85_77),.res(r85_78),.clk(clk),.wout(w85_78));
	PE pe85_79(.x(x79),.w(w85_78),.acc(r85_78),.res(r85_79),.clk(clk),.wout(w85_79));
	PE pe85_80(.x(x80),.w(w85_79),.acc(r85_79),.res(r85_80),.clk(clk),.wout(w85_80));
	PE pe85_81(.x(x81),.w(w85_80),.acc(r85_80),.res(r85_81),.clk(clk),.wout(w85_81));
	PE pe85_82(.x(x82),.w(w85_81),.acc(r85_81),.res(r85_82),.clk(clk),.wout(w85_82));
	PE pe85_83(.x(x83),.w(w85_82),.acc(r85_82),.res(r85_83),.clk(clk),.wout(w85_83));
	PE pe85_84(.x(x84),.w(w85_83),.acc(r85_83),.res(r85_84),.clk(clk),.wout(w85_84));
	PE pe85_85(.x(x85),.w(w85_84),.acc(r85_84),.res(r85_85),.clk(clk),.wout(w85_85));
	PE pe85_86(.x(x86),.w(w85_85),.acc(r85_85),.res(r85_86),.clk(clk),.wout(w85_86));
	PE pe85_87(.x(x87),.w(w85_86),.acc(r85_86),.res(r85_87),.clk(clk),.wout(w85_87));
	PE pe85_88(.x(x88),.w(w85_87),.acc(r85_87),.res(r85_88),.clk(clk),.wout(w85_88));
	PE pe85_89(.x(x89),.w(w85_88),.acc(r85_88),.res(r85_89),.clk(clk),.wout(w85_89));
	PE pe85_90(.x(x90),.w(w85_89),.acc(r85_89),.res(r85_90),.clk(clk),.wout(w85_90));
	PE pe85_91(.x(x91),.w(w85_90),.acc(r85_90),.res(r85_91),.clk(clk),.wout(w85_91));
	PE pe85_92(.x(x92),.w(w85_91),.acc(r85_91),.res(r85_92),.clk(clk),.wout(w85_92));
	PE pe85_93(.x(x93),.w(w85_92),.acc(r85_92),.res(r85_93),.clk(clk),.wout(w85_93));
	PE pe85_94(.x(x94),.w(w85_93),.acc(r85_93),.res(r85_94),.clk(clk),.wout(w85_94));
	PE pe85_95(.x(x95),.w(w85_94),.acc(r85_94),.res(r85_95),.clk(clk),.wout(w85_95));
	PE pe85_96(.x(x96),.w(w85_95),.acc(r85_95),.res(r85_96),.clk(clk),.wout(w85_96));
	PE pe85_97(.x(x97),.w(w85_96),.acc(r85_96),.res(r85_97),.clk(clk),.wout(w85_97));
	PE pe85_98(.x(x98),.w(w85_97),.acc(r85_97),.res(r85_98),.clk(clk),.wout(w85_98));
	PE pe85_99(.x(x99),.w(w85_98),.acc(r85_98),.res(r85_99),.clk(clk),.wout(w85_99));
	PE pe85_100(.x(x100),.w(w85_99),.acc(r85_99),.res(r85_100),.clk(clk),.wout(w85_100));
	PE pe85_101(.x(x101),.w(w85_100),.acc(r85_100),.res(r85_101),.clk(clk),.wout(w85_101));
	PE pe85_102(.x(x102),.w(w85_101),.acc(r85_101),.res(r85_102),.clk(clk),.wout(w85_102));
	PE pe85_103(.x(x103),.w(w85_102),.acc(r85_102),.res(r85_103),.clk(clk),.wout(w85_103));
	PE pe85_104(.x(x104),.w(w85_103),.acc(r85_103),.res(r85_104),.clk(clk),.wout(w85_104));
	PE pe85_105(.x(x105),.w(w85_104),.acc(r85_104),.res(r85_105),.clk(clk),.wout(w85_105));
	PE pe85_106(.x(x106),.w(w85_105),.acc(r85_105),.res(r85_106),.clk(clk),.wout(w85_106));
	PE pe85_107(.x(x107),.w(w85_106),.acc(r85_106),.res(r85_107),.clk(clk),.wout(w85_107));
	PE pe85_108(.x(x108),.w(w85_107),.acc(r85_107),.res(r85_108),.clk(clk),.wout(w85_108));
	PE pe85_109(.x(x109),.w(w85_108),.acc(r85_108),.res(r85_109),.clk(clk),.wout(w85_109));
	PE pe85_110(.x(x110),.w(w85_109),.acc(r85_109),.res(r85_110),.clk(clk),.wout(w85_110));
	PE pe85_111(.x(x111),.w(w85_110),.acc(r85_110),.res(r85_111),.clk(clk),.wout(w85_111));
	PE pe85_112(.x(x112),.w(w85_111),.acc(r85_111),.res(r85_112),.clk(clk),.wout(w85_112));
	PE pe85_113(.x(x113),.w(w85_112),.acc(r85_112),.res(r85_113),.clk(clk),.wout(w85_113));
	PE pe85_114(.x(x114),.w(w85_113),.acc(r85_113),.res(r85_114),.clk(clk),.wout(w85_114));
	PE pe85_115(.x(x115),.w(w85_114),.acc(r85_114),.res(r85_115),.clk(clk),.wout(w85_115));
	PE pe85_116(.x(x116),.w(w85_115),.acc(r85_115),.res(r85_116),.clk(clk),.wout(w85_116));
	PE pe85_117(.x(x117),.w(w85_116),.acc(r85_116),.res(r85_117),.clk(clk),.wout(w85_117));
	PE pe85_118(.x(x118),.w(w85_117),.acc(r85_117),.res(r85_118),.clk(clk),.wout(w85_118));
	PE pe85_119(.x(x119),.w(w85_118),.acc(r85_118),.res(r85_119),.clk(clk),.wout(w85_119));
	PE pe85_120(.x(x120),.w(w85_119),.acc(r85_119),.res(r85_120),.clk(clk),.wout(w85_120));
	PE pe85_121(.x(x121),.w(w85_120),.acc(r85_120),.res(r85_121),.clk(clk),.wout(w85_121));
	PE pe85_122(.x(x122),.w(w85_121),.acc(r85_121),.res(r85_122),.clk(clk),.wout(w85_122));
	PE pe85_123(.x(x123),.w(w85_122),.acc(r85_122),.res(r85_123),.clk(clk),.wout(w85_123));
	PE pe85_124(.x(x124),.w(w85_123),.acc(r85_123),.res(r85_124),.clk(clk),.wout(w85_124));
	PE pe85_125(.x(x125),.w(w85_124),.acc(r85_124),.res(r85_125),.clk(clk),.wout(w85_125));
	PE pe85_126(.x(x126),.w(w85_125),.acc(r85_125),.res(r85_126),.clk(clk),.wout(w85_126));
	PE pe85_127(.x(x127),.w(w85_126),.acc(r85_126),.res(result85),.clk(clk),.wout(weight85));

	PE pe86_0(.x(x0),.w(w86),.acc(32'h0),.res(r86_0),.clk(clk),.wout(w86_0));
	PE pe86_1(.x(x1),.w(w86_0),.acc(r86_0),.res(r86_1),.clk(clk),.wout(w86_1));
	PE pe86_2(.x(x2),.w(w86_1),.acc(r86_1),.res(r86_2),.clk(clk),.wout(w86_2));
	PE pe86_3(.x(x3),.w(w86_2),.acc(r86_2),.res(r86_3),.clk(clk),.wout(w86_3));
	PE pe86_4(.x(x4),.w(w86_3),.acc(r86_3),.res(r86_4),.clk(clk),.wout(w86_4));
	PE pe86_5(.x(x5),.w(w86_4),.acc(r86_4),.res(r86_5),.clk(clk),.wout(w86_5));
	PE pe86_6(.x(x6),.w(w86_5),.acc(r86_5),.res(r86_6),.clk(clk),.wout(w86_6));
	PE pe86_7(.x(x7),.w(w86_6),.acc(r86_6),.res(r86_7),.clk(clk),.wout(w86_7));
	PE pe86_8(.x(x8),.w(w86_7),.acc(r86_7),.res(r86_8),.clk(clk),.wout(w86_8));
	PE pe86_9(.x(x9),.w(w86_8),.acc(r86_8),.res(r86_9),.clk(clk),.wout(w86_9));
	PE pe86_10(.x(x10),.w(w86_9),.acc(r86_9),.res(r86_10),.clk(clk),.wout(w86_10));
	PE pe86_11(.x(x11),.w(w86_10),.acc(r86_10),.res(r86_11),.clk(clk),.wout(w86_11));
	PE pe86_12(.x(x12),.w(w86_11),.acc(r86_11),.res(r86_12),.clk(clk),.wout(w86_12));
	PE pe86_13(.x(x13),.w(w86_12),.acc(r86_12),.res(r86_13),.clk(clk),.wout(w86_13));
	PE pe86_14(.x(x14),.w(w86_13),.acc(r86_13),.res(r86_14),.clk(clk),.wout(w86_14));
	PE pe86_15(.x(x15),.w(w86_14),.acc(r86_14),.res(r86_15),.clk(clk),.wout(w86_15));
	PE pe86_16(.x(x16),.w(w86_15),.acc(r86_15),.res(r86_16),.clk(clk),.wout(w86_16));
	PE pe86_17(.x(x17),.w(w86_16),.acc(r86_16),.res(r86_17),.clk(clk),.wout(w86_17));
	PE pe86_18(.x(x18),.w(w86_17),.acc(r86_17),.res(r86_18),.clk(clk),.wout(w86_18));
	PE pe86_19(.x(x19),.w(w86_18),.acc(r86_18),.res(r86_19),.clk(clk),.wout(w86_19));
	PE pe86_20(.x(x20),.w(w86_19),.acc(r86_19),.res(r86_20),.clk(clk),.wout(w86_20));
	PE pe86_21(.x(x21),.w(w86_20),.acc(r86_20),.res(r86_21),.clk(clk),.wout(w86_21));
	PE pe86_22(.x(x22),.w(w86_21),.acc(r86_21),.res(r86_22),.clk(clk),.wout(w86_22));
	PE pe86_23(.x(x23),.w(w86_22),.acc(r86_22),.res(r86_23),.clk(clk),.wout(w86_23));
	PE pe86_24(.x(x24),.w(w86_23),.acc(r86_23),.res(r86_24),.clk(clk),.wout(w86_24));
	PE pe86_25(.x(x25),.w(w86_24),.acc(r86_24),.res(r86_25),.clk(clk),.wout(w86_25));
	PE pe86_26(.x(x26),.w(w86_25),.acc(r86_25),.res(r86_26),.clk(clk),.wout(w86_26));
	PE pe86_27(.x(x27),.w(w86_26),.acc(r86_26),.res(r86_27),.clk(clk),.wout(w86_27));
	PE pe86_28(.x(x28),.w(w86_27),.acc(r86_27),.res(r86_28),.clk(clk),.wout(w86_28));
	PE pe86_29(.x(x29),.w(w86_28),.acc(r86_28),.res(r86_29),.clk(clk),.wout(w86_29));
	PE pe86_30(.x(x30),.w(w86_29),.acc(r86_29),.res(r86_30),.clk(clk),.wout(w86_30));
	PE pe86_31(.x(x31),.w(w86_30),.acc(r86_30),.res(r86_31),.clk(clk),.wout(w86_31));
	PE pe86_32(.x(x32),.w(w86_31),.acc(r86_31),.res(r86_32),.clk(clk),.wout(w86_32));
	PE pe86_33(.x(x33),.w(w86_32),.acc(r86_32),.res(r86_33),.clk(clk),.wout(w86_33));
	PE pe86_34(.x(x34),.w(w86_33),.acc(r86_33),.res(r86_34),.clk(clk),.wout(w86_34));
	PE pe86_35(.x(x35),.w(w86_34),.acc(r86_34),.res(r86_35),.clk(clk),.wout(w86_35));
	PE pe86_36(.x(x36),.w(w86_35),.acc(r86_35),.res(r86_36),.clk(clk),.wout(w86_36));
	PE pe86_37(.x(x37),.w(w86_36),.acc(r86_36),.res(r86_37),.clk(clk),.wout(w86_37));
	PE pe86_38(.x(x38),.w(w86_37),.acc(r86_37),.res(r86_38),.clk(clk),.wout(w86_38));
	PE pe86_39(.x(x39),.w(w86_38),.acc(r86_38),.res(r86_39),.clk(clk),.wout(w86_39));
	PE pe86_40(.x(x40),.w(w86_39),.acc(r86_39),.res(r86_40),.clk(clk),.wout(w86_40));
	PE pe86_41(.x(x41),.w(w86_40),.acc(r86_40),.res(r86_41),.clk(clk),.wout(w86_41));
	PE pe86_42(.x(x42),.w(w86_41),.acc(r86_41),.res(r86_42),.clk(clk),.wout(w86_42));
	PE pe86_43(.x(x43),.w(w86_42),.acc(r86_42),.res(r86_43),.clk(clk),.wout(w86_43));
	PE pe86_44(.x(x44),.w(w86_43),.acc(r86_43),.res(r86_44),.clk(clk),.wout(w86_44));
	PE pe86_45(.x(x45),.w(w86_44),.acc(r86_44),.res(r86_45),.clk(clk),.wout(w86_45));
	PE pe86_46(.x(x46),.w(w86_45),.acc(r86_45),.res(r86_46),.clk(clk),.wout(w86_46));
	PE pe86_47(.x(x47),.w(w86_46),.acc(r86_46),.res(r86_47),.clk(clk),.wout(w86_47));
	PE pe86_48(.x(x48),.w(w86_47),.acc(r86_47),.res(r86_48),.clk(clk),.wout(w86_48));
	PE pe86_49(.x(x49),.w(w86_48),.acc(r86_48),.res(r86_49),.clk(clk),.wout(w86_49));
	PE pe86_50(.x(x50),.w(w86_49),.acc(r86_49),.res(r86_50),.clk(clk),.wout(w86_50));
	PE pe86_51(.x(x51),.w(w86_50),.acc(r86_50),.res(r86_51),.clk(clk),.wout(w86_51));
	PE pe86_52(.x(x52),.w(w86_51),.acc(r86_51),.res(r86_52),.clk(clk),.wout(w86_52));
	PE pe86_53(.x(x53),.w(w86_52),.acc(r86_52),.res(r86_53),.clk(clk),.wout(w86_53));
	PE pe86_54(.x(x54),.w(w86_53),.acc(r86_53),.res(r86_54),.clk(clk),.wout(w86_54));
	PE pe86_55(.x(x55),.w(w86_54),.acc(r86_54),.res(r86_55),.clk(clk),.wout(w86_55));
	PE pe86_56(.x(x56),.w(w86_55),.acc(r86_55),.res(r86_56),.clk(clk),.wout(w86_56));
	PE pe86_57(.x(x57),.w(w86_56),.acc(r86_56),.res(r86_57),.clk(clk),.wout(w86_57));
	PE pe86_58(.x(x58),.w(w86_57),.acc(r86_57),.res(r86_58),.clk(clk),.wout(w86_58));
	PE pe86_59(.x(x59),.w(w86_58),.acc(r86_58),.res(r86_59),.clk(clk),.wout(w86_59));
	PE pe86_60(.x(x60),.w(w86_59),.acc(r86_59),.res(r86_60),.clk(clk),.wout(w86_60));
	PE pe86_61(.x(x61),.w(w86_60),.acc(r86_60),.res(r86_61),.clk(clk),.wout(w86_61));
	PE pe86_62(.x(x62),.w(w86_61),.acc(r86_61),.res(r86_62),.clk(clk),.wout(w86_62));
	PE pe86_63(.x(x63),.w(w86_62),.acc(r86_62),.res(r86_63),.clk(clk),.wout(w86_63));
	PE pe86_64(.x(x64),.w(w86_63),.acc(r86_63),.res(r86_64),.clk(clk),.wout(w86_64));
	PE pe86_65(.x(x65),.w(w86_64),.acc(r86_64),.res(r86_65),.clk(clk),.wout(w86_65));
	PE pe86_66(.x(x66),.w(w86_65),.acc(r86_65),.res(r86_66),.clk(clk),.wout(w86_66));
	PE pe86_67(.x(x67),.w(w86_66),.acc(r86_66),.res(r86_67),.clk(clk),.wout(w86_67));
	PE pe86_68(.x(x68),.w(w86_67),.acc(r86_67),.res(r86_68),.clk(clk),.wout(w86_68));
	PE pe86_69(.x(x69),.w(w86_68),.acc(r86_68),.res(r86_69),.clk(clk),.wout(w86_69));
	PE pe86_70(.x(x70),.w(w86_69),.acc(r86_69),.res(r86_70),.clk(clk),.wout(w86_70));
	PE pe86_71(.x(x71),.w(w86_70),.acc(r86_70),.res(r86_71),.clk(clk),.wout(w86_71));
	PE pe86_72(.x(x72),.w(w86_71),.acc(r86_71),.res(r86_72),.clk(clk),.wout(w86_72));
	PE pe86_73(.x(x73),.w(w86_72),.acc(r86_72),.res(r86_73),.clk(clk),.wout(w86_73));
	PE pe86_74(.x(x74),.w(w86_73),.acc(r86_73),.res(r86_74),.clk(clk),.wout(w86_74));
	PE pe86_75(.x(x75),.w(w86_74),.acc(r86_74),.res(r86_75),.clk(clk),.wout(w86_75));
	PE pe86_76(.x(x76),.w(w86_75),.acc(r86_75),.res(r86_76),.clk(clk),.wout(w86_76));
	PE pe86_77(.x(x77),.w(w86_76),.acc(r86_76),.res(r86_77),.clk(clk),.wout(w86_77));
	PE pe86_78(.x(x78),.w(w86_77),.acc(r86_77),.res(r86_78),.clk(clk),.wout(w86_78));
	PE pe86_79(.x(x79),.w(w86_78),.acc(r86_78),.res(r86_79),.clk(clk),.wout(w86_79));
	PE pe86_80(.x(x80),.w(w86_79),.acc(r86_79),.res(r86_80),.clk(clk),.wout(w86_80));
	PE pe86_81(.x(x81),.w(w86_80),.acc(r86_80),.res(r86_81),.clk(clk),.wout(w86_81));
	PE pe86_82(.x(x82),.w(w86_81),.acc(r86_81),.res(r86_82),.clk(clk),.wout(w86_82));
	PE pe86_83(.x(x83),.w(w86_82),.acc(r86_82),.res(r86_83),.clk(clk),.wout(w86_83));
	PE pe86_84(.x(x84),.w(w86_83),.acc(r86_83),.res(r86_84),.clk(clk),.wout(w86_84));
	PE pe86_85(.x(x85),.w(w86_84),.acc(r86_84),.res(r86_85),.clk(clk),.wout(w86_85));
	PE pe86_86(.x(x86),.w(w86_85),.acc(r86_85),.res(r86_86),.clk(clk),.wout(w86_86));
	PE pe86_87(.x(x87),.w(w86_86),.acc(r86_86),.res(r86_87),.clk(clk),.wout(w86_87));
	PE pe86_88(.x(x88),.w(w86_87),.acc(r86_87),.res(r86_88),.clk(clk),.wout(w86_88));
	PE pe86_89(.x(x89),.w(w86_88),.acc(r86_88),.res(r86_89),.clk(clk),.wout(w86_89));
	PE pe86_90(.x(x90),.w(w86_89),.acc(r86_89),.res(r86_90),.clk(clk),.wout(w86_90));
	PE pe86_91(.x(x91),.w(w86_90),.acc(r86_90),.res(r86_91),.clk(clk),.wout(w86_91));
	PE pe86_92(.x(x92),.w(w86_91),.acc(r86_91),.res(r86_92),.clk(clk),.wout(w86_92));
	PE pe86_93(.x(x93),.w(w86_92),.acc(r86_92),.res(r86_93),.clk(clk),.wout(w86_93));
	PE pe86_94(.x(x94),.w(w86_93),.acc(r86_93),.res(r86_94),.clk(clk),.wout(w86_94));
	PE pe86_95(.x(x95),.w(w86_94),.acc(r86_94),.res(r86_95),.clk(clk),.wout(w86_95));
	PE pe86_96(.x(x96),.w(w86_95),.acc(r86_95),.res(r86_96),.clk(clk),.wout(w86_96));
	PE pe86_97(.x(x97),.w(w86_96),.acc(r86_96),.res(r86_97),.clk(clk),.wout(w86_97));
	PE pe86_98(.x(x98),.w(w86_97),.acc(r86_97),.res(r86_98),.clk(clk),.wout(w86_98));
	PE pe86_99(.x(x99),.w(w86_98),.acc(r86_98),.res(r86_99),.clk(clk),.wout(w86_99));
	PE pe86_100(.x(x100),.w(w86_99),.acc(r86_99),.res(r86_100),.clk(clk),.wout(w86_100));
	PE pe86_101(.x(x101),.w(w86_100),.acc(r86_100),.res(r86_101),.clk(clk),.wout(w86_101));
	PE pe86_102(.x(x102),.w(w86_101),.acc(r86_101),.res(r86_102),.clk(clk),.wout(w86_102));
	PE pe86_103(.x(x103),.w(w86_102),.acc(r86_102),.res(r86_103),.clk(clk),.wout(w86_103));
	PE pe86_104(.x(x104),.w(w86_103),.acc(r86_103),.res(r86_104),.clk(clk),.wout(w86_104));
	PE pe86_105(.x(x105),.w(w86_104),.acc(r86_104),.res(r86_105),.clk(clk),.wout(w86_105));
	PE pe86_106(.x(x106),.w(w86_105),.acc(r86_105),.res(r86_106),.clk(clk),.wout(w86_106));
	PE pe86_107(.x(x107),.w(w86_106),.acc(r86_106),.res(r86_107),.clk(clk),.wout(w86_107));
	PE pe86_108(.x(x108),.w(w86_107),.acc(r86_107),.res(r86_108),.clk(clk),.wout(w86_108));
	PE pe86_109(.x(x109),.w(w86_108),.acc(r86_108),.res(r86_109),.clk(clk),.wout(w86_109));
	PE pe86_110(.x(x110),.w(w86_109),.acc(r86_109),.res(r86_110),.clk(clk),.wout(w86_110));
	PE pe86_111(.x(x111),.w(w86_110),.acc(r86_110),.res(r86_111),.clk(clk),.wout(w86_111));
	PE pe86_112(.x(x112),.w(w86_111),.acc(r86_111),.res(r86_112),.clk(clk),.wout(w86_112));
	PE pe86_113(.x(x113),.w(w86_112),.acc(r86_112),.res(r86_113),.clk(clk),.wout(w86_113));
	PE pe86_114(.x(x114),.w(w86_113),.acc(r86_113),.res(r86_114),.clk(clk),.wout(w86_114));
	PE pe86_115(.x(x115),.w(w86_114),.acc(r86_114),.res(r86_115),.clk(clk),.wout(w86_115));
	PE pe86_116(.x(x116),.w(w86_115),.acc(r86_115),.res(r86_116),.clk(clk),.wout(w86_116));
	PE pe86_117(.x(x117),.w(w86_116),.acc(r86_116),.res(r86_117),.clk(clk),.wout(w86_117));
	PE pe86_118(.x(x118),.w(w86_117),.acc(r86_117),.res(r86_118),.clk(clk),.wout(w86_118));
	PE pe86_119(.x(x119),.w(w86_118),.acc(r86_118),.res(r86_119),.clk(clk),.wout(w86_119));
	PE pe86_120(.x(x120),.w(w86_119),.acc(r86_119),.res(r86_120),.clk(clk),.wout(w86_120));
	PE pe86_121(.x(x121),.w(w86_120),.acc(r86_120),.res(r86_121),.clk(clk),.wout(w86_121));
	PE pe86_122(.x(x122),.w(w86_121),.acc(r86_121),.res(r86_122),.clk(clk),.wout(w86_122));
	PE pe86_123(.x(x123),.w(w86_122),.acc(r86_122),.res(r86_123),.clk(clk),.wout(w86_123));
	PE pe86_124(.x(x124),.w(w86_123),.acc(r86_123),.res(r86_124),.clk(clk),.wout(w86_124));
	PE pe86_125(.x(x125),.w(w86_124),.acc(r86_124),.res(r86_125),.clk(clk),.wout(w86_125));
	PE pe86_126(.x(x126),.w(w86_125),.acc(r86_125),.res(r86_126),.clk(clk),.wout(w86_126));
	PE pe86_127(.x(x127),.w(w86_126),.acc(r86_126),.res(result86),.clk(clk),.wout(weight86));

	PE pe87_0(.x(x0),.w(w87),.acc(32'h0),.res(r87_0),.clk(clk),.wout(w87_0));
	PE pe87_1(.x(x1),.w(w87_0),.acc(r87_0),.res(r87_1),.clk(clk),.wout(w87_1));
	PE pe87_2(.x(x2),.w(w87_1),.acc(r87_1),.res(r87_2),.clk(clk),.wout(w87_2));
	PE pe87_3(.x(x3),.w(w87_2),.acc(r87_2),.res(r87_3),.clk(clk),.wout(w87_3));
	PE pe87_4(.x(x4),.w(w87_3),.acc(r87_3),.res(r87_4),.clk(clk),.wout(w87_4));
	PE pe87_5(.x(x5),.w(w87_4),.acc(r87_4),.res(r87_5),.clk(clk),.wout(w87_5));
	PE pe87_6(.x(x6),.w(w87_5),.acc(r87_5),.res(r87_6),.clk(clk),.wout(w87_6));
	PE pe87_7(.x(x7),.w(w87_6),.acc(r87_6),.res(r87_7),.clk(clk),.wout(w87_7));
	PE pe87_8(.x(x8),.w(w87_7),.acc(r87_7),.res(r87_8),.clk(clk),.wout(w87_8));
	PE pe87_9(.x(x9),.w(w87_8),.acc(r87_8),.res(r87_9),.clk(clk),.wout(w87_9));
	PE pe87_10(.x(x10),.w(w87_9),.acc(r87_9),.res(r87_10),.clk(clk),.wout(w87_10));
	PE pe87_11(.x(x11),.w(w87_10),.acc(r87_10),.res(r87_11),.clk(clk),.wout(w87_11));
	PE pe87_12(.x(x12),.w(w87_11),.acc(r87_11),.res(r87_12),.clk(clk),.wout(w87_12));
	PE pe87_13(.x(x13),.w(w87_12),.acc(r87_12),.res(r87_13),.clk(clk),.wout(w87_13));
	PE pe87_14(.x(x14),.w(w87_13),.acc(r87_13),.res(r87_14),.clk(clk),.wout(w87_14));
	PE pe87_15(.x(x15),.w(w87_14),.acc(r87_14),.res(r87_15),.clk(clk),.wout(w87_15));
	PE pe87_16(.x(x16),.w(w87_15),.acc(r87_15),.res(r87_16),.clk(clk),.wout(w87_16));
	PE pe87_17(.x(x17),.w(w87_16),.acc(r87_16),.res(r87_17),.clk(clk),.wout(w87_17));
	PE pe87_18(.x(x18),.w(w87_17),.acc(r87_17),.res(r87_18),.clk(clk),.wout(w87_18));
	PE pe87_19(.x(x19),.w(w87_18),.acc(r87_18),.res(r87_19),.clk(clk),.wout(w87_19));
	PE pe87_20(.x(x20),.w(w87_19),.acc(r87_19),.res(r87_20),.clk(clk),.wout(w87_20));
	PE pe87_21(.x(x21),.w(w87_20),.acc(r87_20),.res(r87_21),.clk(clk),.wout(w87_21));
	PE pe87_22(.x(x22),.w(w87_21),.acc(r87_21),.res(r87_22),.clk(clk),.wout(w87_22));
	PE pe87_23(.x(x23),.w(w87_22),.acc(r87_22),.res(r87_23),.clk(clk),.wout(w87_23));
	PE pe87_24(.x(x24),.w(w87_23),.acc(r87_23),.res(r87_24),.clk(clk),.wout(w87_24));
	PE pe87_25(.x(x25),.w(w87_24),.acc(r87_24),.res(r87_25),.clk(clk),.wout(w87_25));
	PE pe87_26(.x(x26),.w(w87_25),.acc(r87_25),.res(r87_26),.clk(clk),.wout(w87_26));
	PE pe87_27(.x(x27),.w(w87_26),.acc(r87_26),.res(r87_27),.clk(clk),.wout(w87_27));
	PE pe87_28(.x(x28),.w(w87_27),.acc(r87_27),.res(r87_28),.clk(clk),.wout(w87_28));
	PE pe87_29(.x(x29),.w(w87_28),.acc(r87_28),.res(r87_29),.clk(clk),.wout(w87_29));
	PE pe87_30(.x(x30),.w(w87_29),.acc(r87_29),.res(r87_30),.clk(clk),.wout(w87_30));
	PE pe87_31(.x(x31),.w(w87_30),.acc(r87_30),.res(r87_31),.clk(clk),.wout(w87_31));
	PE pe87_32(.x(x32),.w(w87_31),.acc(r87_31),.res(r87_32),.clk(clk),.wout(w87_32));
	PE pe87_33(.x(x33),.w(w87_32),.acc(r87_32),.res(r87_33),.clk(clk),.wout(w87_33));
	PE pe87_34(.x(x34),.w(w87_33),.acc(r87_33),.res(r87_34),.clk(clk),.wout(w87_34));
	PE pe87_35(.x(x35),.w(w87_34),.acc(r87_34),.res(r87_35),.clk(clk),.wout(w87_35));
	PE pe87_36(.x(x36),.w(w87_35),.acc(r87_35),.res(r87_36),.clk(clk),.wout(w87_36));
	PE pe87_37(.x(x37),.w(w87_36),.acc(r87_36),.res(r87_37),.clk(clk),.wout(w87_37));
	PE pe87_38(.x(x38),.w(w87_37),.acc(r87_37),.res(r87_38),.clk(clk),.wout(w87_38));
	PE pe87_39(.x(x39),.w(w87_38),.acc(r87_38),.res(r87_39),.clk(clk),.wout(w87_39));
	PE pe87_40(.x(x40),.w(w87_39),.acc(r87_39),.res(r87_40),.clk(clk),.wout(w87_40));
	PE pe87_41(.x(x41),.w(w87_40),.acc(r87_40),.res(r87_41),.clk(clk),.wout(w87_41));
	PE pe87_42(.x(x42),.w(w87_41),.acc(r87_41),.res(r87_42),.clk(clk),.wout(w87_42));
	PE pe87_43(.x(x43),.w(w87_42),.acc(r87_42),.res(r87_43),.clk(clk),.wout(w87_43));
	PE pe87_44(.x(x44),.w(w87_43),.acc(r87_43),.res(r87_44),.clk(clk),.wout(w87_44));
	PE pe87_45(.x(x45),.w(w87_44),.acc(r87_44),.res(r87_45),.clk(clk),.wout(w87_45));
	PE pe87_46(.x(x46),.w(w87_45),.acc(r87_45),.res(r87_46),.clk(clk),.wout(w87_46));
	PE pe87_47(.x(x47),.w(w87_46),.acc(r87_46),.res(r87_47),.clk(clk),.wout(w87_47));
	PE pe87_48(.x(x48),.w(w87_47),.acc(r87_47),.res(r87_48),.clk(clk),.wout(w87_48));
	PE pe87_49(.x(x49),.w(w87_48),.acc(r87_48),.res(r87_49),.clk(clk),.wout(w87_49));
	PE pe87_50(.x(x50),.w(w87_49),.acc(r87_49),.res(r87_50),.clk(clk),.wout(w87_50));
	PE pe87_51(.x(x51),.w(w87_50),.acc(r87_50),.res(r87_51),.clk(clk),.wout(w87_51));
	PE pe87_52(.x(x52),.w(w87_51),.acc(r87_51),.res(r87_52),.clk(clk),.wout(w87_52));
	PE pe87_53(.x(x53),.w(w87_52),.acc(r87_52),.res(r87_53),.clk(clk),.wout(w87_53));
	PE pe87_54(.x(x54),.w(w87_53),.acc(r87_53),.res(r87_54),.clk(clk),.wout(w87_54));
	PE pe87_55(.x(x55),.w(w87_54),.acc(r87_54),.res(r87_55),.clk(clk),.wout(w87_55));
	PE pe87_56(.x(x56),.w(w87_55),.acc(r87_55),.res(r87_56),.clk(clk),.wout(w87_56));
	PE pe87_57(.x(x57),.w(w87_56),.acc(r87_56),.res(r87_57),.clk(clk),.wout(w87_57));
	PE pe87_58(.x(x58),.w(w87_57),.acc(r87_57),.res(r87_58),.clk(clk),.wout(w87_58));
	PE pe87_59(.x(x59),.w(w87_58),.acc(r87_58),.res(r87_59),.clk(clk),.wout(w87_59));
	PE pe87_60(.x(x60),.w(w87_59),.acc(r87_59),.res(r87_60),.clk(clk),.wout(w87_60));
	PE pe87_61(.x(x61),.w(w87_60),.acc(r87_60),.res(r87_61),.clk(clk),.wout(w87_61));
	PE pe87_62(.x(x62),.w(w87_61),.acc(r87_61),.res(r87_62),.clk(clk),.wout(w87_62));
	PE pe87_63(.x(x63),.w(w87_62),.acc(r87_62),.res(r87_63),.clk(clk),.wout(w87_63));
	PE pe87_64(.x(x64),.w(w87_63),.acc(r87_63),.res(r87_64),.clk(clk),.wout(w87_64));
	PE pe87_65(.x(x65),.w(w87_64),.acc(r87_64),.res(r87_65),.clk(clk),.wout(w87_65));
	PE pe87_66(.x(x66),.w(w87_65),.acc(r87_65),.res(r87_66),.clk(clk),.wout(w87_66));
	PE pe87_67(.x(x67),.w(w87_66),.acc(r87_66),.res(r87_67),.clk(clk),.wout(w87_67));
	PE pe87_68(.x(x68),.w(w87_67),.acc(r87_67),.res(r87_68),.clk(clk),.wout(w87_68));
	PE pe87_69(.x(x69),.w(w87_68),.acc(r87_68),.res(r87_69),.clk(clk),.wout(w87_69));
	PE pe87_70(.x(x70),.w(w87_69),.acc(r87_69),.res(r87_70),.clk(clk),.wout(w87_70));
	PE pe87_71(.x(x71),.w(w87_70),.acc(r87_70),.res(r87_71),.clk(clk),.wout(w87_71));
	PE pe87_72(.x(x72),.w(w87_71),.acc(r87_71),.res(r87_72),.clk(clk),.wout(w87_72));
	PE pe87_73(.x(x73),.w(w87_72),.acc(r87_72),.res(r87_73),.clk(clk),.wout(w87_73));
	PE pe87_74(.x(x74),.w(w87_73),.acc(r87_73),.res(r87_74),.clk(clk),.wout(w87_74));
	PE pe87_75(.x(x75),.w(w87_74),.acc(r87_74),.res(r87_75),.clk(clk),.wout(w87_75));
	PE pe87_76(.x(x76),.w(w87_75),.acc(r87_75),.res(r87_76),.clk(clk),.wout(w87_76));
	PE pe87_77(.x(x77),.w(w87_76),.acc(r87_76),.res(r87_77),.clk(clk),.wout(w87_77));
	PE pe87_78(.x(x78),.w(w87_77),.acc(r87_77),.res(r87_78),.clk(clk),.wout(w87_78));
	PE pe87_79(.x(x79),.w(w87_78),.acc(r87_78),.res(r87_79),.clk(clk),.wout(w87_79));
	PE pe87_80(.x(x80),.w(w87_79),.acc(r87_79),.res(r87_80),.clk(clk),.wout(w87_80));
	PE pe87_81(.x(x81),.w(w87_80),.acc(r87_80),.res(r87_81),.clk(clk),.wout(w87_81));
	PE pe87_82(.x(x82),.w(w87_81),.acc(r87_81),.res(r87_82),.clk(clk),.wout(w87_82));
	PE pe87_83(.x(x83),.w(w87_82),.acc(r87_82),.res(r87_83),.clk(clk),.wout(w87_83));
	PE pe87_84(.x(x84),.w(w87_83),.acc(r87_83),.res(r87_84),.clk(clk),.wout(w87_84));
	PE pe87_85(.x(x85),.w(w87_84),.acc(r87_84),.res(r87_85),.clk(clk),.wout(w87_85));
	PE pe87_86(.x(x86),.w(w87_85),.acc(r87_85),.res(r87_86),.clk(clk),.wout(w87_86));
	PE pe87_87(.x(x87),.w(w87_86),.acc(r87_86),.res(r87_87),.clk(clk),.wout(w87_87));
	PE pe87_88(.x(x88),.w(w87_87),.acc(r87_87),.res(r87_88),.clk(clk),.wout(w87_88));
	PE pe87_89(.x(x89),.w(w87_88),.acc(r87_88),.res(r87_89),.clk(clk),.wout(w87_89));
	PE pe87_90(.x(x90),.w(w87_89),.acc(r87_89),.res(r87_90),.clk(clk),.wout(w87_90));
	PE pe87_91(.x(x91),.w(w87_90),.acc(r87_90),.res(r87_91),.clk(clk),.wout(w87_91));
	PE pe87_92(.x(x92),.w(w87_91),.acc(r87_91),.res(r87_92),.clk(clk),.wout(w87_92));
	PE pe87_93(.x(x93),.w(w87_92),.acc(r87_92),.res(r87_93),.clk(clk),.wout(w87_93));
	PE pe87_94(.x(x94),.w(w87_93),.acc(r87_93),.res(r87_94),.clk(clk),.wout(w87_94));
	PE pe87_95(.x(x95),.w(w87_94),.acc(r87_94),.res(r87_95),.clk(clk),.wout(w87_95));
	PE pe87_96(.x(x96),.w(w87_95),.acc(r87_95),.res(r87_96),.clk(clk),.wout(w87_96));
	PE pe87_97(.x(x97),.w(w87_96),.acc(r87_96),.res(r87_97),.clk(clk),.wout(w87_97));
	PE pe87_98(.x(x98),.w(w87_97),.acc(r87_97),.res(r87_98),.clk(clk),.wout(w87_98));
	PE pe87_99(.x(x99),.w(w87_98),.acc(r87_98),.res(r87_99),.clk(clk),.wout(w87_99));
	PE pe87_100(.x(x100),.w(w87_99),.acc(r87_99),.res(r87_100),.clk(clk),.wout(w87_100));
	PE pe87_101(.x(x101),.w(w87_100),.acc(r87_100),.res(r87_101),.clk(clk),.wout(w87_101));
	PE pe87_102(.x(x102),.w(w87_101),.acc(r87_101),.res(r87_102),.clk(clk),.wout(w87_102));
	PE pe87_103(.x(x103),.w(w87_102),.acc(r87_102),.res(r87_103),.clk(clk),.wout(w87_103));
	PE pe87_104(.x(x104),.w(w87_103),.acc(r87_103),.res(r87_104),.clk(clk),.wout(w87_104));
	PE pe87_105(.x(x105),.w(w87_104),.acc(r87_104),.res(r87_105),.clk(clk),.wout(w87_105));
	PE pe87_106(.x(x106),.w(w87_105),.acc(r87_105),.res(r87_106),.clk(clk),.wout(w87_106));
	PE pe87_107(.x(x107),.w(w87_106),.acc(r87_106),.res(r87_107),.clk(clk),.wout(w87_107));
	PE pe87_108(.x(x108),.w(w87_107),.acc(r87_107),.res(r87_108),.clk(clk),.wout(w87_108));
	PE pe87_109(.x(x109),.w(w87_108),.acc(r87_108),.res(r87_109),.clk(clk),.wout(w87_109));
	PE pe87_110(.x(x110),.w(w87_109),.acc(r87_109),.res(r87_110),.clk(clk),.wout(w87_110));
	PE pe87_111(.x(x111),.w(w87_110),.acc(r87_110),.res(r87_111),.clk(clk),.wout(w87_111));
	PE pe87_112(.x(x112),.w(w87_111),.acc(r87_111),.res(r87_112),.clk(clk),.wout(w87_112));
	PE pe87_113(.x(x113),.w(w87_112),.acc(r87_112),.res(r87_113),.clk(clk),.wout(w87_113));
	PE pe87_114(.x(x114),.w(w87_113),.acc(r87_113),.res(r87_114),.clk(clk),.wout(w87_114));
	PE pe87_115(.x(x115),.w(w87_114),.acc(r87_114),.res(r87_115),.clk(clk),.wout(w87_115));
	PE pe87_116(.x(x116),.w(w87_115),.acc(r87_115),.res(r87_116),.clk(clk),.wout(w87_116));
	PE pe87_117(.x(x117),.w(w87_116),.acc(r87_116),.res(r87_117),.clk(clk),.wout(w87_117));
	PE pe87_118(.x(x118),.w(w87_117),.acc(r87_117),.res(r87_118),.clk(clk),.wout(w87_118));
	PE pe87_119(.x(x119),.w(w87_118),.acc(r87_118),.res(r87_119),.clk(clk),.wout(w87_119));
	PE pe87_120(.x(x120),.w(w87_119),.acc(r87_119),.res(r87_120),.clk(clk),.wout(w87_120));
	PE pe87_121(.x(x121),.w(w87_120),.acc(r87_120),.res(r87_121),.clk(clk),.wout(w87_121));
	PE pe87_122(.x(x122),.w(w87_121),.acc(r87_121),.res(r87_122),.clk(clk),.wout(w87_122));
	PE pe87_123(.x(x123),.w(w87_122),.acc(r87_122),.res(r87_123),.clk(clk),.wout(w87_123));
	PE pe87_124(.x(x124),.w(w87_123),.acc(r87_123),.res(r87_124),.clk(clk),.wout(w87_124));
	PE pe87_125(.x(x125),.w(w87_124),.acc(r87_124),.res(r87_125),.clk(clk),.wout(w87_125));
	PE pe87_126(.x(x126),.w(w87_125),.acc(r87_125),.res(r87_126),.clk(clk),.wout(w87_126));
	PE pe87_127(.x(x127),.w(w87_126),.acc(r87_126),.res(result87),.clk(clk),.wout(weight87));

	PE pe88_0(.x(x0),.w(w88),.acc(32'h0),.res(r88_0),.clk(clk),.wout(w88_0));
	PE pe88_1(.x(x1),.w(w88_0),.acc(r88_0),.res(r88_1),.clk(clk),.wout(w88_1));
	PE pe88_2(.x(x2),.w(w88_1),.acc(r88_1),.res(r88_2),.clk(clk),.wout(w88_2));
	PE pe88_3(.x(x3),.w(w88_2),.acc(r88_2),.res(r88_3),.clk(clk),.wout(w88_3));
	PE pe88_4(.x(x4),.w(w88_3),.acc(r88_3),.res(r88_4),.clk(clk),.wout(w88_4));
	PE pe88_5(.x(x5),.w(w88_4),.acc(r88_4),.res(r88_5),.clk(clk),.wout(w88_5));
	PE pe88_6(.x(x6),.w(w88_5),.acc(r88_5),.res(r88_6),.clk(clk),.wout(w88_6));
	PE pe88_7(.x(x7),.w(w88_6),.acc(r88_6),.res(r88_7),.clk(clk),.wout(w88_7));
	PE pe88_8(.x(x8),.w(w88_7),.acc(r88_7),.res(r88_8),.clk(clk),.wout(w88_8));
	PE pe88_9(.x(x9),.w(w88_8),.acc(r88_8),.res(r88_9),.clk(clk),.wout(w88_9));
	PE pe88_10(.x(x10),.w(w88_9),.acc(r88_9),.res(r88_10),.clk(clk),.wout(w88_10));
	PE pe88_11(.x(x11),.w(w88_10),.acc(r88_10),.res(r88_11),.clk(clk),.wout(w88_11));
	PE pe88_12(.x(x12),.w(w88_11),.acc(r88_11),.res(r88_12),.clk(clk),.wout(w88_12));
	PE pe88_13(.x(x13),.w(w88_12),.acc(r88_12),.res(r88_13),.clk(clk),.wout(w88_13));
	PE pe88_14(.x(x14),.w(w88_13),.acc(r88_13),.res(r88_14),.clk(clk),.wout(w88_14));
	PE pe88_15(.x(x15),.w(w88_14),.acc(r88_14),.res(r88_15),.clk(clk),.wout(w88_15));
	PE pe88_16(.x(x16),.w(w88_15),.acc(r88_15),.res(r88_16),.clk(clk),.wout(w88_16));
	PE pe88_17(.x(x17),.w(w88_16),.acc(r88_16),.res(r88_17),.clk(clk),.wout(w88_17));
	PE pe88_18(.x(x18),.w(w88_17),.acc(r88_17),.res(r88_18),.clk(clk),.wout(w88_18));
	PE pe88_19(.x(x19),.w(w88_18),.acc(r88_18),.res(r88_19),.clk(clk),.wout(w88_19));
	PE pe88_20(.x(x20),.w(w88_19),.acc(r88_19),.res(r88_20),.clk(clk),.wout(w88_20));
	PE pe88_21(.x(x21),.w(w88_20),.acc(r88_20),.res(r88_21),.clk(clk),.wout(w88_21));
	PE pe88_22(.x(x22),.w(w88_21),.acc(r88_21),.res(r88_22),.clk(clk),.wout(w88_22));
	PE pe88_23(.x(x23),.w(w88_22),.acc(r88_22),.res(r88_23),.clk(clk),.wout(w88_23));
	PE pe88_24(.x(x24),.w(w88_23),.acc(r88_23),.res(r88_24),.clk(clk),.wout(w88_24));
	PE pe88_25(.x(x25),.w(w88_24),.acc(r88_24),.res(r88_25),.clk(clk),.wout(w88_25));
	PE pe88_26(.x(x26),.w(w88_25),.acc(r88_25),.res(r88_26),.clk(clk),.wout(w88_26));
	PE pe88_27(.x(x27),.w(w88_26),.acc(r88_26),.res(r88_27),.clk(clk),.wout(w88_27));
	PE pe88_28(.x(x28),.w(w88_27),.acc(r88_27),.res(r88_28),.clk(clk),.wout(w88_28));
	PE pe88_29(.x(x29),.w(w88_28),.acc(r88_28),.res(r88_29),.clk(clk),.wout(w88_29));
	PE pe88_30(.x(x30),.w(w88_29),.acc(r88_29),.res(r88_30),.clk(clk),.wout(w88_30));
	PE pe88_31(.x(x31),.w(w88_30),.acc(r88_30),.res(r88_31),.clk(clk),.wout(w88_31));
	PE pe88_32(.x(x32),.w(w88_31),.acc(r88_31),.res(r88_32),.clk(clk),.wout(w88_32));
	PE pe88_33(.x(x33),.w(w88_32),.acc(r88_32),.res(r88_33),.clk(clk),.wout(w88_33));
	PE pe88_34(.x(x34),.w(w88_33),.acc(r88_33),.res(r88_34),.clk(clk),.wout(w88_34));
	PE pe88_35(.x(x35),.w(w88_34),.acc(r88_34),.res(r88_35),.clk(clk),.wout(w88_35));
	PE pe88_36(.x(x36),.w(w88_35),.acc(r88_35),.res(r88_36),.clk(clk),.wout(w88_36));
	PE pe88_37(.x(x37),.w(w88_36),.acc(r88_36),.res(r88_37),.clk(clk),.wout(w88_37));
	PE pe88_38(.x(x38),.w(w88_37),.acc(r88_37),.res(r88_38),.clk(clk),.wout(w88_38));
	PE pe88_39(.x(x39),.w(w88_38),.acc(r88_38),.res(r88_39),.clk(clk),.wout(w88_39));
	PE pe88_40(.x(x40),.w(w88_39),.acc(r88_39),.res(r88_40),.clk(clk),.wout(w88_40));
	PE pe88_41(.x(x41),.w(w88_40),.acc(r88_40),.res(r88_41),.clk(clk),.wout(w88_41));
	PE pe88_42(.x(x42),.w(w88_41),.acc(r88_41),.res(r88_42),.clk(clk),.wout(w88_42));
	PE pe88_43(.x(x43),.w(w88_42),.acc(r88_42),.res(r88_43),.clk(clk),.wout(w88_43));
	PE pe88_44(.x(x44),.w(w88_43),.acc(r88_43),.res(r88_44),.clk(clk),.wout(w88_44));
	PE pe88_45(.x(x45),.w(w88_44),.acc(r88_44),.res(r88_45),.clk(clk),.wout(w88_45));
	PE pe88_46(.x(x46),.w(w88_45),.acc(r88_45),.res(r88_46),.clk(clk),.wout(w88_46));
	PE pe88_47(.x(x47),.w(w88_46),.acc(r88_46),.res(r88_47),.clk(clk),.wout(w88_47));
	PE pe88_48(.x(x48),.w(w88_47),.acc(r88_47),.res(r88_48),.clk(clk),.wout(w88_48));
	PE pe88_49(.x(x49),.w(w88_48),.acc(r88_48),.res(r88_49),.clk(clk),.wout(w88_49));
	PE pe88_50(.x(x50),.w(w88_49),.acc(r88_49),.res(r88_50),.clk(clk),.wout(w88_50));
	PE pe88_51(.x(x51),.w(w88_50),.acc(r88_50),.res(r88_51),.clk(clk),.wout(w88_51));
	PE pe88_52(.x(x52),.w(w88_51),.acc(r88_51),.res(r88_52),.clk(clk),.wout(w88_52));
	PE pe88_53(.x(x53),.w(w88_52),.acc(r88_52),.res(r88_53),.clk(clk),.wout(w88_53));
	PE pe88_54(.x(x54),.w(w88_53),.acc(r88_53),.res(r88_54),.clk(clk),.wout(w88_54));
	PE pe88_55(.x(x55),.w(w88_54),.acc(r88_54),.res(r88_55),.clk(clk),.wout(w88_55));
	PE pe88_56(.x(x56),.w(w88_55),.acc(r88_55),.res(r88_56),.clk(clk),.wout(w88_56));
	PE pe88_57(.x(x57),.w(w88_56),.acc(r88_56),.res(r88_57),.clk(clk),.wout(w88_57));
	PE pe88_58(.x(x58),.w(w88_57),.acc(r88_57),.res(r88_58),.clk(clk),.wout(w88_58));
	PE pe88_59(.x(x59),.w(w88_58),.acc(r88_58),.res(r88_59),.clk(clk),.wout(w88_59));
	PE pe88_60(.x(x60),.w(w88_59),.acc(r88_59),.res(r88_60),.clk(clk),.wout(w88_60));
	PE pe88_61(.x(x61),.w(w88_60),.acc(r88_60),.res(r88_61),.clk(clk),.wout(w88_61));
	PE pe88_62(.x(x62),.w(w88_61),.acc(r88_61),.res(r88_62),.clk(clk),.wout(w88_62));
	PE pe88_63(.x(x63),.w(w88_62),.acc(r88_62),.res(r88_63),.clk(clk),.wout(w88_63));
	PE pe88_64(.x(x64),.w(w88_63),.acc(r88_63),.res(r88_64),.clk(clk),.wout(w88_64));
	PE pe88_65(.x(x65),.w(w88_64),.acc(r88_64),.res(r88_65),.clk(clk),.wout(w88_65));
	PE pe88_66(.x(x66),.w(w88_65),.acc(r88_65),.res(r88_66),.clk(clk),.wout(w88_66));
	PE pe88_67(.x(x67),.w(w88_66),.acc(r88_66),.res(r88_67),.clk(clk),.wout(w88_67));
	PE pe88_68(.x(x68),.w(w88_67),.acc(r88_67),.res(r88_68),.clk(clk),.wout(w88_68));
	PE pe88_69(.x(x69),.w(w88_68),.acc(r88_68),.res(r88_69),.clk(clk),.wout(w88_69));
	PE pe88_70(.x(x70),.w(w88_69),.acc(r88_69),.res(r88_70),.clk(clk),.wout(w88_70));
	PE pe88_71(.x(x71),.w(w88_70),.acc(r88_70),.res(r88_71),.clk(clk),.wout(w88_71));
	PE pe88_72(.x(x72),.w(w88_71),.acc(r88_71),.res(r88_72),.clk(clk),.wout(w88_72));
	PE pe88_73(.x(x73),.w(w88_72),.acc(r88_72),.res(r88_73),.clk(clk),.wout(w88_73));
	PE pe88_74(.x(x74),.w(w88_73),.acc(r88_73),.res(r88_74),.clk(clk),.wout(w88_74));
	PE pe88_75(.x(x75),.w(w88_74),.acc(r88_74),.res(r88_75),.clk(clk),.wout(w88_75));
	PE pe88_76(.x(x76),.w(w88_75),.acc(r88_75),.res(r88_76),.clk(clk),.wout(w88_76));
	PE pe88_77(.x(x77),.w(w88_76),.acc(r88_76),.res(r88_77),.clk(clk),.wout(w88_77));
	PE pe88_78(.x(x78),.w(w88_77),.acc(r88_77),.res(r88_78),.clk(clk),.wout(w88_78));
	PE pe88_79(.x(x79),.w(w88_78),.acc(r88_78),.res(r88_79),.clk(clk),.wout(w88_79));
	PE pe88_80(.x(x80),.w(w88_79),.acc(r88_79),.res(r88_80),.clk(clk),.wout(w88_80));
	PE pe88_81(.x(x81),.w(w88_80),.acc(r88_80),.res(r88_81),.clk(clk),.wout(w88_81));
	PE pe88_82(.x(x82),.w(w88_81),.acc(r88_81),.res(r88_82),.clk(clk),.wout(w88_82));
	PE pe88_83(.x(x83),.w(w88_82),.acc(r88_82),.res(r88_83),.clk(clk),.wout(w88_83));
	PE pe88_84(.x(x84),.w(w88_83),.acc(r88_83),.res(r88_84),.clk(clk),.wout(w88_84));
	PE pe88_85(.x(x85),.w(w88_84),.acc(r88_84),.res(r88_85),.clk(clk),.wout(w88_85));
	PE pe88_86(.x(x86),.w(w88_85),.acc(r88_85),.res(r88_86),.clk(clk),.wout(w88_86));
	PE pe88_87(.x(x87),.w(w88_86),.acc(r88_86),.res(r88_87),.clk(clk),.wout(w88_87));
	PE pe88_88(.x(x88),.w(w88_87),.acc(r88_87),.res(r88_88),.clk(clk),.wout(w88_88));
	PE pe88_89(.x(x89),.w(w88_88),.acc(r88_88),.res(r88_89),.clk(clk),.wout(w88_89));
	PE pe88_90(.x(x90),.w(w88_89),.acc(r88_89),.res(r88_90),.clk(clk),.wout(w88_90));
	PE pe88_91(.x(x91),.w(w88_90),.acc(r88_90),.res(r88_91),.clk(clk),.wout(w88_91));
	PE pe88_92(.x(x92),.w(w88_91),.acc(r88_91),.res(r88_92),.clk(clk),.wout(w88_92));
	PE pe88_93(.x(x93),.w(w88_92),.acc(r88_92),.res(r88_93),.clk(clk),.wout(w88_93));
	PE pe88_94(.x(x94),.w(w88_93),.acc(r88_93),.res(r88_94),.clk(clk),.wout(w88_94));
	PE pe88_95(.x(x95),.w(w88_94),.acc(r88_94),.res(r88_95),.clk(clk),.wout(w88_95));
	PE pe88_96(.x(x96),.w(w88_95),.acc(r88_95),.res(r88_96),.clk(clk),.wout(w88_96));
	PE pe88_97(.x(x97),.w(w88_96),.acc(r88_96),.res(r88_97),.clk(clk),.wout(w88_97));
	PE pe88_98(.x(x98),.w(w88_97),.acc(r88_97),.res(r88_98),.clk(clk),.wout(w88_98));
	PE pe88_99(.x(x99),.w(w88_98),.acc(r88_98),.res(r88_99),.clk(clk),.wout(w88_99));
	PE pe88_100(.x(x100),.w(w88_99),.acc(r88_99),.res(r88_100),.clk(clk),.wout(w88_100));
	PE pe88_101(.x(x101),.w(w88_100),.acc(r88_100),.res(r88_101),.clk(clk),.wout(w88_101));
	PE pe88_102(.x(x102),.w(w88_101),.acc(r88_101),.res(r88_102),.clk(clk),.wout(w88_102));
	PE pe88_103(.x(x103),.w(w88_102),.acc(r88_102),.res(r88_103),.clk(clk),.wout(w88_103));
	PE pe88_104(.x(x104),.w(w88_103),.acc(r88_103),.res(r88_104),.clk(clk),.wout(w88_104));
	PE pe88_105(.x(x105),.w(w88_104),.acc(r88_104),.res(r88_105),.clk(clk),.wout(w88_105));
	PE pe88_106(.x(x106),.w(w88_105),.acc(r88_105),.res(r88_106),.clk(clk),.wout(w88_106));
	PE pe88_107(.x(x107),.w(w88_106),.acc(r88_106),.res(r88_107),.clk(clk),.wout(w88_107));
	PE pe88_108(.x(x108),.w(w88_107),.acc(r88_107),.res(r88_108),.clk(clk),.wout(w88_108));
	PE pe88_109(.x(x109),.w(w88_108),.acc(r88_108),.res(r88_109),.clk(clk),.wout(w88_109));
	PE pe88_110(.x(x110),.w(w88_109),.acc(r88_109),.res(r88_110),.clk(clk),.wout(w88_110));
	PE pe88_111(.x(x111),.w(w88_110),.acc(r88_110),.res(r88_111),.clk(clk),.wout(w88_111));
	PE pe88_112(.x(x112),.w(w88_111),.acc(r88_111),.res(r88_112),.clk(clk),.wout(w88_112));
	PE pe88_113(.x(x113),.w(w88_112),.acc(r88_112),.res(r88_113),.clk(clk),.wout(w88_113));
	PE pe88_114(.x(x114),.w(w88_113),.acc(r88_113),.res(r88_114),.clk(clk),.wout(w88_114));
	PE pe88_115(.x(x115),.w(w88_114),.acc(r88_114),.res(r88_115),.clk(clk),.wout(w88_115));
	PE pe88_116(.x(x116),.w(w88_115),.acc(r88_115),.res(r88_116),.clk(clk),.wout(w88_116));
	PE pe88_117(.x(x117),.w(w88_116),.acc(r88_116),.res(r88_117),.clk(clk),.wout(w88_117));
	PE pe88_118(.x(x118),.w(w88_117),.acc(r88_117),.res(r88_118),.clk(clk),.wout(w88_118));
	PE pe88_119(.x(x119),.w(w88_118),.acc(r88_118),.res(r88_119),.clk(clk),.wout(w88_119));
	PE pe88_120(.x(x120),.w(w88_119),.acc(r88_119),.res(r88_120),.clk(clk),.wout(w88_120));
	PE pe88_121(.x(x121),.w(w88_120),.acc(r88_120),.res(r88_121),.clk(clk),.wout(w88_121));
	PE pe88_122(.x(x122),.w(w88_121),.acc(r88_121),.res(r88_122),.clk(clk),.wout(w88_122));
	PE pe88_123(.x(x123),.w(w88_122),.acc(r88_122),.res(r88_123),.clk(clk),.wout(w88_123));
	PE pe88_124(.x(x124),.w(w88_123),.acc(r88_123),.res(r88_124),.clk(clk),.wout(w88_124));
	PE pe88_125(.x(x125),.w(w88_124),.acc(r88_124),.res(r88_125),.clk(clk),.wout(w88_125));
	PE pe88_126(.x(x126),.w(w88_125),.acc(r88_125),.res(r88_126),.clk(clk),.wout(w88_126));
	PE pe88_127(.x(x127),.w(w88_126),.acc(r88_126),.res(result88),.clk(clk),.wout(weight88));

	PE pe89_0(.x(x0),.w(w89),.acc(32'h0),.res(r89_0),.clk(clk),.wout(w89_0));
	PE pe89_1(.x(x1),.w(w89_0),.acc(r89_0),.res(r89_1),.clk(clk),.wout(w89_1));
	PE pe89_2(.x(x2),.w(w89_1),.acc(r89_1),.res(r89_2),.clk(clk),.wout(w89_2));
	PE pe89_3(.x(x3),.w(w89_2),.acc(r89_2),.res(r89_3),.clk(clk),.wout(w89_3));
	PE pe89_4(.x(x4),.w(w89_3),.acc(r89_3),.res(r89_4),.clk(clk),.wout(w89_4));
	PE pe89_5(.x(x5),.w(w89_4),.acc(r89_4),.res(r89_5),.clk(clk),.wout(w89_5));
	PE pe89_6(.x(x6),.w(w89_5),.acc(r89_5),.res(r89_6),.clk(clk),.wout(w89_6));
	PE pe89_7(.x(x7),.w(w89_6),.acc(r89_6),.res(r89_7),.clk(clk),.wout(w89_7));
	PE pe89_8(.x(x8),.w(w89_7),.acc(r89_7),.res(r89_8),.clk(clk),.wout(w89_8));
	PE pe89_9(.x(x9),.w(w89_8),.acc(r89_8),.res(r89_9),.clk(clk),.wout(w89_9));
	PE pe89_10(.x(x10),.w(w89_9),.acc(r89_9),.res(r89_10),.clk(clk),.wout(w89_10));
	PE pe89_11(.x(x11),.w(w89_10),.acc(r89_10),.res(r89_11),.clk(clk),.wout(w89_11));
	PE pe89_12(.x(x12),.w(w89_11),.acc(r89_11),.res(r89_12),.clk(clk),.wout(w89_12));
	PE pe89_13(.x(x13),.w(w89_12),.acc(r89_12),.res(r89_13),.clk(clk),.wout(w89_13));
	PE pe89_14(.x(x14),.w(w89_13),.acc(r89_13),.res(r89_14),.clk(clk),.wout(w89_14));
	PE pe89_15(.x(x15),.w(w89_14),.acc(r89_14),.res(r89_15),.clk(clk),.wout(w89_15));
	PE pe89_16(.x(x16),.w(w89_15),.acc(r89_15),.res(r89_16),.clk(clk),.wout(w89_16));
	PE pe89_17(.x(x17),.w(w89_16),.acc(r89_16),.res(r89_17),.clk(clk),.wout(w89_17));
	PE pe89_18(.x(x18),.w(w89_17),.acc(r89_17),.res(r89_18),.clk(clk),.wout(w89_18));
	PE pe89_19(.x(x19),.w(w89_18),.acc(r89_18),.res(r89_19),.clk(clk),.wout(w89_19));
	PE pe89_20(.x(x20),.w(w89_19),.acc(r89_19),.res(r89_20),.clk(clk),.wout(w89_20));
	PE pe89_21(.x(x21),.w(w89_20),.acc(r89_20),.res(r89_21),.clk(clk),.wout(w89_21));
	PE pe89_22(.x(x22),.w(w89_21),.acc(r89_21),.res(r89_22),.clk(clk),.wout(w89_22));
	PE pe89_23(.x(x23),.w(w89_22),.acc(r89_22),.res(r89_23),.clk(clk),.wout(w89_23));
	PE pe89_24(.x(x24),.w(w89_23),.acc(r89_23),.res(r89_24),.clk(clk),.wout(w89_24));
	PE pe89_25(.x(x25),.w(w89_24),.acc(r89_24),.res(r89_25),.clk(clk),.wout(w89_25));
	PE pe89_26(.x(x26),.w(w89_25),.acc(r89_25),.res(r89_26),.clk(clk),.wout(w89_26));
	PE pe89_27(.x(x27),.w(w89_26),.acc(r89_26),.res(r89_27),.clk(clk),.wout(w89_27));
	PE pe89_28(.x(x28),.w(w89_27),.acc(r89_27),.res(r89_28),.clk(clk),.wout(w89_28));
	PE pe89_29(.x(x29),.w(w89_28),.acc(r89_28),.res(r89_29),.clk(clk),.wout(w89_29));
	PE pe89_30(.x(x30),.w(w89_29),.acc(r89_29),.res(r89_30),.clk(clk),.wout(w89_30));
	PE pe89_31(.x(x31),.w(w89_30),.acc(r89_30),.res(r89_31),.clk(clk),.wout(w89_31));
	PE pe89_32(.x(x32),.w(w89_31),.acc(r89_31),.res(r89_32),.clk(clk),.wout(w89_32));
	PE pe89_33(.x(x33),.w(w89_32),.acc(r89_32),.res(r89_33),.clk(clk),.wout(w89_33));
	PE pe89_34(.x(x34),.w(w89_33),.acc(r89_33),.res(r89_34),.clk(clk),.wout(w89_34));
	PE pe89_35(.x(x35),.w(w89_34),.acc(r89_34),.res(r89_35),.clk(clk),.wout(w89_35));
	PE pe89_36(.x(x36),.w(w89_35),.acc(r89_35),.res(r89_36),.clk(clk),.wout(w89_36));
	PE pe89_37(.x(x37),.w(w89_36),.acc(r89_36),.res(r89_37),.clk(clk),.wout(w89_37));
	PE pe89_38(.x(x38),.w(w89_37),.acc(r89_37),.res(r89_38),.clk(clk),.wout(w89_38));
	PE pe89_39(.x(x39),.w(w89_38),.acc(r89_38),.res(r89_39),.clk(clk),.wout(w89_39));
	PE pe89_40(.x(x40),.w(w89_39),.acc(r89_39),.res(r89_40),.clk(clk),.wout(w89_40));
	PE pe89_41(.x(x41),.w(w89_40),.acc(r89_40),.res(r89_41),.clk(clk),.wout(w89_41));
	PE pe89_42(.x(x42),.w(w89_41),.acc(r89_41),.res(r89_42),.clk(clk),.wout(w89_42));
	PE pe89_43(.x(x43),.w(w89_42),.acc(r89_42),.res(r89_43),.clk(clk),.wout(w89_43));
	PE pe89_44(.x(x44),.w(w89_43),.acc(r89_43),.res(r89_44),.clk(clk),.wout(w89_44));
	PE pe89_45(.x(x45),.w(w89_44),.acc(r89_44),.res(r89_45),.clk(clk),.wout(w89_45));
	PE pe89_46(.x(x46),.w(w89_45),.acc(r89_45),.res(r89_46),.clk(clk),.wout(w89_46));
	PE pe89_47(.x(x47),.w(w89_46),.acc(r89_46),.res(r89_47),.clk(clk),.wout(w89_47));
	PE pe89_48(.x(x48),.w(w89_47),.acc(r89_47),.res(r89_48),.clk(clk),.wout(w89_48));
	PE pe89_49(.x(x49),.w(w89_48),.acc(r89_48),.res(r89_49),.clk(clk),.wout(w89_49));
	PE pe89_50(.x(x50),.w(w89_49),.acc(r89_49),.res(r89_50),.clk(clk),.wout(w89_50));
	PE pe89_51(.x(x51),.w(w89_50),.acc(r89_50),.res(r89_51),.clk(clk),.wout(w89_51));
	PE pe89_52(.x(x52),.w(w89_51),.acc(r89_51),.res(r89_52),.clk(clk),.wout(w89_52));
	PE pe89_53(.x(x53),.w(w89_52),.acc(r89_52),.res(r89_53),.clk(clk),.wout(w89_53));
	PE pe89_54(.x(x54),.w(w89_53),.acc(r89_53),.res(r89_54),.clk(clk),.wout(w89_54));
	PE pe89_55(.x(x55),.w(w89_54),.acc(r89_54),.res(r89_55),.clk(clk),.wout(w89_55));
	PE pe89_56(.x(x56),.w(w89_55),.acc(r89_55),.res(r89_56),.clk(clk),.wout(w89_56));
	PE pe89_57(.x(x57),.w(w89_56),.acc(r89_56),.res(r89_57),.clk(clk),.wout(w89_57));
	PE pe89_58(.x(x58),.w(w89_57),.acc(r89_57),.res(r89_58),.clk(clk),.wout(w89_58));
	PE pe89_59(.x(x59),.w(w89_58),.acc(r89_58),.res(r89_59),.clk(clk),.wout(w89_59));
	PE pe89_60(.x(x60),.w(w89_59),.acc(r89_59),.res(r89_60),.clk(clk),.wout(w89_60));
	PE pe89_61(.x(x61),.w(w89_60),.acc(r89_60),.res(r89_61),.clk(clk),.wout(w89_61));
	PE pe89_62(.x(x62),.w(w89_61),.acc(r89_61),.res(r89_62),.clk(clk),.wout(w89_62));
	PE pe89_63(.x(x63),.w(w89_62),.acc(r89_62),.res(r89_63),.clk(clk),.wout(w89_63));
	PE pe89_64(.x(x64),.w(w89_63),.acc(r89_63),.res(r89_64),.clk(clk),.wout(w89_64));
	PE pe89_65(.x(x65),.w(w89_64),.acc(r89_64),.res(r89_65),.clk(clk),.wout(w89_65));
	PE pe89_66(.x(x66),.w(w89_65),.acc(r89_65),.res(r89_66),.clk(clk),.wout(w89_66));
	PE pe89_67(.x(x67),.w(w89_66),.acc(r89_66),.res(r89_67),.clk(clk),.wout(w89_67));
	PE pe89_68(.x(x68),.w(w89_67),.acc(r89_67),.res(r89_68),.clk(clk),.wout(w89_68));
	PE pe89_69(.x(x69),.w(w89_68),.acc(r89_68),.res(r89_69),.clk(clk),.wout(w89_69));
	PE pe89_70(.x(x70),.w(w89_69),.acc(r89_69),.res(r89_70),.clk(clk),.wout(w89_70));
	PE pe89_71(.x(x71),.w(w89_70),.acc(r89_70),.res(r89_71),.clk(clk),.wout(w89_71));
	PE pe89_72(.x(x72),.w(w89_71),.acc(r89_71),.res(r89_72),.clk(clk),.wout(w89_72));
	PE pe89_73(.x(x73),.w(w89_72),.acc(r89_72),.res(r89_73),.clk(clk),.wout(w89_73));
	PE pe89_74(.x(x74),.w(w89_73),.acc(r89_73),.res(r89_74),.clk(clk),.wout(w89_74));
	PE pe89_75(.x(x75),.w(w89_74),.acc(r89_74),.res(r89_75),.clk(clk),.wout(w89_75));
	PE pe89_76(.x(x76),.w(w89_75),.acc(r89_75),.res(r89_76),.clk(clk),.wout(w89_76));
	PE pe89_77(.x(x77),.w(w89_76),.acc(r89_76),.res(r89_77),.clk(clk),.wout(w89_77));
	PE pe89_78(.x(x78),.w(w89_77),.acc(r89_77),.res(r89_78),.clk(clk),.wout(w89_78));
	PE pe89_79(.x(x79),.w(w89_78),.acc(r89_78),.res(r89_79),.clk(clk),.wout(w89_79));
	PE pe89_80(.x(x80),.w(w89_79),.acc(r89_79),.res(r89_80),.clk(clk),.wout(w89_80));
	PE pe89_81(.x(x81),.w(w89_80),.acc(r89_80),.res(r89_81),.clk(clk),.wout(w89_81));
	PE pe89_82(.x(x82),.w(w89_81),.acc(r89_81),.res(r89_82),.clk(clk),.wout(w89_82));
	PE pe89_83(.x(x83),.w(w89_82),.acc(r89_82),.res(r89_83),.clk(clk),.wout(w89_83));
	PE pe89_84(.x(x84),.w(w89_83),.acc(r89_83),.res(r89_84),.clk(clk),.wout(w89_84));
	PE pe89_85(.x(x85),.w(w89_84),.acc(r89_84),.res(r89_85),.clk(clk),.wout(w89_85));
	PE pe89_86(.x(x86),.w(w89_85),.acc(r89_85),.res(r89_86),.clk(clk),.wout(w89_86));
	PE pe89_87(.x(x87),.w(w89_86),.acc(r89_86),.res(r89_87),.clk(clk),.wout(w89_87));
	PE pe89_88(.x(x88),.w(w89_87),.acc(r89_87),.res(r89_88),.clk(clk),.wout(w89_88));
	PE pe89_89(.x(x89),.w(w89_88),.acc(r89_88),.res(r89_89),.clk(clk),.wout(w89_89));
	PE pe89_90(.x(x90),.w(w89_89),.acc(r89_89),.res(r89_90),.clk(clk),.wout(w89_90));
	PE pe89_91(.x(x91),.w(w89_90),.acc(r89_90),.res(r89_91),.clk(clk),.wout(w89_91));
	PE pe89_92(.x(x92),.w(w89_91),.acc(r89_91),.res(r89_92),.clk(clk),.wout(w89_92));
	PE pe89_93(.x(x93),.w(w89_92),.acc(r89_92),.res(r89_93),.clk(clk),.wout(w89_93));
	PE pe89_94(.x(x94),.w(w89_93),.acc(r89_93),.res(r89_94),.clk(clk),.wout(w89_94));
	PE pe89_95(.x(x95),.w(w89_94),.acc(r89_94),.res(r89_95),.clk(clk),.wout(w89_95));
	PE pe89_96(.x(x96),.w(w89_95),.acc(r89_95),.res(r89_96),.clk(clk),.wout(w89_96));
	PE pe89_97(.x(x97),.w(w89_96),.acc(r89_96),.res(r89_97),.clk(clk),.wout(w89_97));
	PE pe89_98(.x(x98),.w(w89_97),.acc(r89_97),.res(r89_98),.clk(clk),.wout(w89_98));
	PE pe89_99(.x(x99),.w(w89_98),.acc(r89_98),.res(r89_99),.clk(clk),.wout(w89_99));
	PE pe89_100(.x(x100),.w(w89_99),.acc(r89_99),.res(r89_100),.clk(clk),.wout(w89_100));
	PE pe89_101(.x(x101),.w(w89_100),.acc(r89_100),.res(r89_101),.clk(clk),.wout(w89_101));
	PE pe89_102(.x(x102),.w(w89_101),.acc(r89_101),.res(r89_102),.clk(clk),.wout(w89_102));
	PE pe89_103(.x(x103),.w(w89_102),.acc(r89_102),.res(r89_103),.clk(clk),.wout(w89_103));
	PE pe89_104(.x(x104),.w(w89_103),.acc(r89_103),.res(r89_104),.clk(clk),.wout(w89_104));
	PE pe89_105(.x(x105),.w(w89_104),.acc(r89_104),.res(r89_105),.clk(clk),.wout(w89_105));
	PE pe89_106(.x(x106),.w(w89_105),.acc(r89_105),.res(r89_106),.clk(clk),.wout(w89_106));
	PE pe89_107(.x(x107),.w(w89_106),.acc(r89_106),.res(r89_107),.clk(clk),.wout(w89_107));
	PE pe89_108(.x(x108),.w(w89_107),.acc(r89_107),.res(r89_108),.clk(clk),.wout(w89_108));
	PE pe89_109(.x(x109),.w(w89_108),.acc(r89_108),.res(r89_109),.clk(clk),.wout(w89_109));
	PE pe89_110(.x(x110),.w(w89_109),.acc(r89_109),.res(r89_110),.clk(clk),.wout(w89_110));
	PE pe89_111(.x(x111),.w(w89_110),.acc(r89_110),.res(r89_111),.clk(clk),.wout(w89_111));
	PE pe89_112(.x(x112),.w(w89_111),.acc(r89_111),.res(r89_112),.clk(clk),.wout(w89_112));
	PE pe89_113(.x(x113),.w(w89_112),.acc(r89_112),.res(r89_113),.clk(clk),.wout(w89_113));
	PE pe89_114(.x(x114),.w(w89_113),.acc(r89_113),.res(r89_114),.clk(clk),.wout(w89_114));
	PE pe89_115(.x(x115),.w(w89_114),.acc(r89_114),.res(r89_115),.clk(clk),.wout(w89_115));
	PE pe89_116(.x(x116),.w(w89_115),.acc(r89_115),.res(r89_116),.clk(clk),.wout(w89_116));
	PE pe89_117(.x(x117),.w(w89_116),.acc(r89_116),.res(r89_117),.clk(clk),.wout(w89_117));
	PE pe89_118(.x(x118),.w(w89_117),.acc(r89_117),.res(r89_118),.clk(clk),.wout(w89_118));
	PE pe89_119(.x(x119),.w(w89_118),.acc(r89_118),.res(r89_119),.clk(clk),.wout(w89_119));
	PE pe89_120(.x(x120),.w(w89_119),.acc(r89_119),.res(r89_120),.clk(clk),.wout(w89_120));
	PE pe89_121(.x(x121),.w(w89_120),.acc(r89_120),.res(r89_121),.clk(clk),.wout(w89_121));
	PE pe89_122(.x(x122),.w(w89_121),.acc(r89_121),.res(r89_122),.clk(clk),.wout(w89_122));
	PE pe89_123(.x(x123),.w(w89_122),.acc(r89_122),.res(r89_123),.clk(clk),.wout(w89_123));
	PE pe89_124(.x(x124),.w(w89_123),.acc(r89_123),.res(r89_124),.clk(clk),.wout(w89_124));
	PE pe89_125(.x(x125),.w(w89_124),.acc(r89_124),.res(r89_125),.clk(clk),.wout(w89_125));
	PE pe89_126(.x(x126),.w(w89_125),.acc(r89_125),.res(r89_126),.clk(clk),.wout(w89_126));
	PE pe89_127(.x(x127),.w(w89_126),.acc(r89_126),.res(result89),.clk(clk),.wout(weight89));

	PE pe90_0(.x(x0),.w(w90),.acc(32'h0),.res(r90_0),.clk(clk),.wout(w90_0));
	PE pe90_1(.x(x1),.w(w90_0),.acc(r90_0),.res(r90_1),.clk(clk),.wout(w90_1));
	PE pe90_2(.x(x2),.w(w90_1),.acc(r90_1),.res(r90_2),.clk(clk),.wout(w90_2));
	PE pe90_3(.x(x3),.w(w90_2),.acc(r90_2),.res(r90_3),.clk(clk),.wout(w90_3));
	PE pe90_4(.x(x4),.w(w90_3),.acc(r90_3),.res(r90_4),.clk(clk),.wout(w90_4));
	PE pe90_5(.x(x5),.w(w90_4),.acc(r90_4),.res(r90_5),.clk(clk),.wout(w90_5));
	PE pe90_6(.x(x6),.w(w90_5),.acc(r90_5),.res(r90_6),.clk(clk),.wout(w90_6));
	PE pe90_7(.x(x7),.w(w90_6),.acc(r90_6),.res(r90_7),.clk(clk),.wout(w90_7));
	PE pe90_8(.x(x8),.w(w90_7),.acc(r90_7),.res(r90_8),.clk(clk),.wout(w90_8));
	PE pe90_9(.x(x9),.w(w90_8),.acc(r90_8),.res(r90_9),.clk(clk),.wout(w90_9));
	PE pe90_10(.x(x10),.w(w90_9),.acc(r90_9),.res(r90_10),.clk(clk),.wout(w90_10));
	PE pe90_11(.x(x11),.w(w90_10),.acc(r90_10),.res(r90_11),.clk(clk),.wout(w90_11));
	PE pe90_12(.x(x12),.w(w90_11),.acc(r90_11),.res(r90_12),.clk(clk),.wout(w90_12));
	PE pe90_13(.x(x13),.w(w90_12),.acc(r90_12),.res(r90_13),.clk(clk),.wout(w90_13));
	PE pe90_14(.x(x14),.w(w90_13),.acc(r90_13),.res(r90_14),.clk(clk),.wout(w90_14));
	PE pe90_15(.x(x15),.w(w90_14),.acc(r90_14),.res(r90_15),.clk(clk),.wout(w90_15));
	PE pe90_16(.x(x16),.w(w90_15),.acc(r90_15),.res(r90_16),.clk(clk),.wout(w90_16));
	PE pe90_17(.x(x17),.w(w90_16),.acc(r90_16),.res(r90_17),.clk(clk),.wout(w90_17));
	PE pe90_18(.x(x18),.w(w90_17),.acc(r90_17),.res(r90_18),.clk(clk),.wout(w90_18));
	PE pe90_19(.x(x19),.w(w90_18),.acc(r90_18),.res(r90_19),.clk(clk),.wout(w90_19));
	PE pe90_20(.x(x20),.w(w90_19),.acc(r90_19),.res(r90_20),.clk(clk),.wout(w90_20));
	PE pe90_21(.x(x21),.w(w90_20),.acc(r90_20),.res(r90_21),.clk(clk),.wout(w90_21));
	PE pe90_22(.x(x22),.w(w90_21),.acc(r90_21),.res(r90_22),.clk(clk),.wout(w90_22));
	PE pe90_23(.x(x23),.w(w90_22),.acc(r90_22),.res(r90_23),.clk(clk),.wout(w90_23));
	PE pe90_24(.x(x24),.w(w90_23),.acc(r90_23),.res(r90_24),.clk(clk),.wout(w90_24));
	PE pe90_25(.x(x25),.w(w90_24),.acc(r90_24),.res(r90_25),.clk(clk),.wout(w90_25));
	PE pe90_26(.x(x26),.w(w90_25),.acc(r90_25),.res(r90_26),.clk(clk),.wout(w90_26));
	PE pe90_27(.x(x27),.w(w90_26),.acc(r90_26),.res(r90_27),.clk(clk),.wout(w90_27));
	PE pe90_28(.x(x28),.w(w90_27),.acc(r90_27),.res(r90_28),.clk(clk),.wout(w90_28));
	PE pe90_29(.x(x29),.w(w90_28),.acc(r90_28),.res(r90_29),.clk(clk),.wout(w90_29));
	PE pe90_30(.x(x30),.w(w90_29),.acc(r90_29),.res(r90_30),.clk(clk),.wout(w90_30));
	PE pe90_31(.x(x31),.w(w90_30),.acc(r90_30),.res(r90_31),.clk(clk),.wout(w90_31));
	PE pe90_32(.x(x32),.w(w90_31),.acc(r90_31),.res(r90_32),.clk(clk),.wout(w90_32));
	PE pe90_33(.x(x33),.w(w90_32),.acc(r90_32),.res(r90_33),.clk(clk),.wout(w90_33));
	PE pe90_34(.x(x34),.w(w90_33),.acc(r90_33),.res(r90_34),.clk(clk),.wout(w90_34));
	PE pe90_35(.x(x35),.w(w90_34),.acc(r90_34),.res(r90_35),.clk(clk),.wout(w90_35));
	PE pe90_36(.x(x36),.w(w90_35),.acc(r90_35),.res(r90_36),.clk(clk),.wout(w90_36));
	PE pe90_37(.x(x37),.w(w90_36),.acc(r90_36),.res(r90_37),.clk(clk),.wout(w90_37));
	PE pe90_38(.x(x38),.w(w90_37),.acc(r90_37),.res(r90_38),.clk(clk),.wout(w90_38));
	PE pe90_39(.x(x39),.w(w90_38),.acc(r90_38),.res(r90_39),.clk(clk),.wout(w90_39));
	PE pe90_40(.x(x40),.w(w90_39),.acc(r90_39),.res(r90_40),.clk(clk),.wout(w90_40));
	PE pe90_41(.x(x41),.w(w90_40),.acc(r90_40),.res(r90_41),.clk(clk),.wout(w90_41));
	PE pe90_42(.x(x42),.w(w90_41),.acc(r90_41),.res(r90_42),.clk(clk),.wout(w90_42));
	PE pe90_43(.x(x43),.w(w90_42),.acc(r90_42),.res(r90_43),.clk(clk),.wout(w90_43));
	PE pe90_44(.x(x44),.w(w90_43),.acc(r90_43),.res(r90_44),.clk(clk),.wout(w90_44));
	PE pe90_45(.x(x45),.w(w90_44),.acc(r90_44),.res(r90_45),.clk(clk),.wout(w90_45));
	PE pe90_46(.x(x46),.w(w90_45),.acc(r90_45),.res(r90_46),.clk(clk),.wout(w90_46));
	PE pe90_47(.x(x47),.w(w90_46),.acc(r90_46),.res(r90_47),.clk(clk),.wout(w90_47));
	PE pe90_48(.x(x48),.w(w90_47),.acc(r90_47),.res(r90_48),.clk(clk),.wout(w90_48));
	PE pe90_49(.x(x49),.w(w90_48),.acc(r90_48),.res(r90_49),.clk(clk),.wout(w90_49));
	PE pe90_50(.x(x50),.w(w90_49),.acc(r90_49),.res(r90_50),.clk(clk),.wout(w90_50));
	PE pe90_51(.x(x51),.w(w90_50),.acc(r90_50),.res(r90_51),.clk(clk),.wout(w90_51));
	PE pe90_52(.x(x52),.w(w90_51),.acc(r90_51),.res(r90_52),.clk(clk),.wout(w90_52));
	PE pe90_53(.x(x53),.w(w90_52),.acc(r90_52),.res(r90_53),.clk(clk),.wout(w90_53));
	PE pe90_54(.x(x54),.w(w90_53),.acc(r90_53),.res(r90_54),.clk(clk),.wout(w90_54));
	PE pe90_55(.x(x55),.w(w90_54),.acc(r90_54),.res(r90_55),.clk(clk),.wout(w90_55));
	PE pe90_56(.x(x56),.w(w90_55),.acc(r90_55),.res(r90_56),.clk(clk),.wout(w90_56));
	PE pe90_57(.x(x57),.w(w90_56),.acc(r90_56),.res(r90_57),.clk(clk),.wout(w90_57));
	PE pe90_58(.x(x58),.w(w90_57),.acc(r90_57),.res(r90_58),.clk(clk),.wout(w90_58));
	PE pe90_59(.x(x59),.w(w90_58),.acc(r90_58),.res(r90_59),.clk(clk),.wout(w90_59));
	PE pe90_60(.x(x60),.w(w90_59),.acc(r90_59),.res(r90_60),.clk(clk),.wout(w90_60));
	PE pe90_61(.x(x61),.w(w90_60),.acc(r90_60),.res(r90_61),.clk(clk),.wout(w90_61));
	PE pe90_62(.x(x62),.w(w90_61),.acc(r90_61),.res(r90_62),.clk(clk),.wout(w90_62));
	PE pe90_63(.x(x63),.w(w90_62),.acc(r90_62),.res(r90_63),.clk(clk),.wout(w90_63));
	PE pe90_64(.x(x64),.w(w90_63),.acc(r90_63),.res(r90_64),.clk(clk),.wout(w90_64));
	PE pe90_65(.x(x65),.w(w90_64),.acc(r90_64),.res(r90_65),.clk(clk),.wout(w90_65));
	PE pe90_66(.x(x66),.w(w90_65),.acc(r90_65),.res(r90_66),.clk(clk),.wout(w90_66));
	PE pe90_67(.x(x67),.w(w90_66),.acc(r90_66),.res(r90_67),.clk(clk),.wout(w90_67));
	PE pe90_68(.x(x68),.w(w90_67),.acc(r90_67),.res(r90_68),.clk(clk),.wout(w90_68));
	PE pe90_69(.x(x69),.w(w90_68),.acc(r90_68),.res(r90_69),.clk(clk),.wout(w90_69));
	PE pe90_70(.x(x70),.w(w90_69),.acc(r90_69),.res(r90_70),.clk(clk),.wout(w90_70));
	PE pe90_71(.x(x71),.w(w90_70),.acc(r90_70),.res(r90_71),.clk(clk),.wout(w90_71));
	PE pe90_72(.x(x72),.w(w90_71),.acc(r90_71),.res(r90_72),.clk(clk),.wout(w90_72));
	PE pe90_73(.x(x73),.w(w90_72),.acc(r90_72),.res(r90_73),.clk(clk),.wout(w90_73));
	PE pe90_74(.x(x74),.w(w90_73),.acc(r90_73),.res(r90_74),.clk(clk),.wout(w90_74));
	PE pe90_75(.x(x75),.w(w90_74),.acc(r90_74),.res(r90_75),.clk(clk),.wout(w90_75));
	PE pe90_76(.x(x76),.w(w90_75),.acc(r90_75),.res(r90_76),.clk(clk),.wout(w90_76));
	PE pe90_77(.x(x77),.w(w90_76),.acc(r90_76),.res(r90_77),.clk(clk),.wout(w90_77));
	PE pe90_78(.x(x78),.w(w90_77),.acc(r90_77),.res(r90_78),.clk(clk),.wout(w90_78));
	PE pe90_79(.x(x79),.w(w90_78),.acc(r90_78),.res(r90_79),.clk(clk),.wout(w90_79));
	PE pe90_80(.x(x80),.w(w90_79),.acc(r90_79),.res(r90_80),.clk(clk),.wout(w90_80));
	PE pe90_81(.x(x81),.w(w90_80),.acc(r90_80),.res(r90_81),.clk(clk),.wout(w90_81));
	PE pe90_82(.x(x82),.w(w90_81),.acc(r90_81),.res(r90_82),.clk(clk),.wout(w90_82));
	PE pe90_83(.x(x83),.w(w90_82),.acc(r90_82),.res(r90_83),.clk(clk),.wout(w90_83));
	PE pe90_84(.x(x84),.w(w90_83),.acc(r90_83),.res(r90_84),.clk(clk),.wout(w90_84));
	PE pe90_85(.x(x85),.w(w90_84),.acc(r90_84),.res(r90_85),.clk(clk),.wout(w90_85));
	PE pe90_86(.x(x86),.w(w90_85),.acc(r90_85),.res(r90_86),.clk(clk),.wout(w90_86));
	PE pe90_87(.x(x87),.w(w90_86),.acc(r90_86),.res(r90_87),.clk(clk),.wout(w90_87));
	PE pe90_88(.x(x88),.w(w90_87),.acc(r90_87),.res(r90_88),.clk(clk),.wout(w90_88));
	PE pe90_89(.x(x89),.w(w90_88),.acc(r90_88),.res(r90_89),.clk(clk),.wout(w90_89));
	PE pe90_90(.x(x90),.w(w90_89),.acc(r90_89),.res(r90_90),.clk(clk),.wout(w90_90));
	PE pe90_91(.x(x91),.w(w90_90),.acc(r90_90),.res(r90_91),.clk(clk),.wout(w90_91));
	PE pe90_92(.x(x92),.w(w90_91),.acc(r90_91),.res(r90_92),.clk(clk),.wout(w90_92));
	PE pe90_93(.x(x93),.w(w90_92),.acc(r90_92),.res(r90_93),.clk(clk),.wout(w90_93));
	PE pe90_94(.x(x94),.w(w90_93),.acc(r90_93),.res(r90_94),.clk(clk),.wout(w90_94));
	PE pe90_95(.x(x95),.w(w90_94),.acc(r90_94),.res(r90_95),.clk(clk),.wout(w90_95));
	PE pe90_96(.x(x96),.w(w90_95),.acc(r90_95),.res(r90_96),.clk(clk),.wout(w90_96));
	PE pe90_97(.x(x97),.w(w90_96),.acc(r90_96),.res(r90_97),.clk(clk),.wout(w90_97));
	PE pe90_98(.x(x98),.w(w90_97),.acc(r90_97),.res(r90_98),.clk(clk),.wout(w90_98));
	PE pe90_99(.x(x99),.w(w90_98),.acc(r90_98),.res(r90_99),.clk(clk),.wout(w90_99));
	PE pe90_100(.x(x100),.w(w90_99),.acc(r90_99),.res(r90_100),.clk(clk),.wout(w90_100));
	PE pe90_101(.x(x101),.w(w90_100),.acc(r90_100),.res(r90_101),.clk(clk),.wout(w90_101));
	PE pe90_102(.x(x102),.w(w90_101),.acc(r90_101),.res(r90_102),.clk(clk),.wout(w90_102));
	PE pe90_103(.x(x103),.w(w90_102),.acc(r90_102),.res(r90_103),.clk(clk),.wout(w90_103));
	PE pe90_104(.x(x104),.w(w90_103),.acc(r90_103),.res(r90_104),.clk(clk),.wout(w90_104));
	PE pe90_105(.x(x105),.w(w90_104),.acc(r90_104),.res(r90_105),.clk(clk),.wout(w90_105));
	PE pe90_106(.x(x106),.w(w90_105),.acc(r90_105),.res(r90_106),.clk(clk),.wout(w90_106));
	PE pe90_107(.x(x107),.w(w90_106),.acc(r90_106),.res(r90_107),.clk(clk),.wout(w90_107));
	PE pe90_108(.x(x108),.w(w90_107),.acc(r90_107),.res(r90_108),.clk(clk),.wout(w90_108));
	PE pe90_109(.x(x109),.w(w90_108),.acc(r90_108),.res(r90_109),.clk(clk),.wout(w90_109));
	PE pe90_110(.x(x110),.w(w90_109),.acc(r90_109),.res(r90_110),.clk(clk),.wout(w90_110));
	PE pe90_111(.x(x111),.w(w90_110),.acc(r90_110),.res(r90_111),.clk(clk),.wout(w90_111));
	PE pe90_112(.x(x112),.w(w90_111),.acc(r90_111),.res(r90_112),.clk(clk),.wout(w90_112));
	PE pe90_113(.x(x113),.w(w90_112),.acc(r90_112),.res(r90_113),.clk(clk),.wout(w90_113));
	PE pe90_114(.x(x114),.w(w90_113),.acc(r90_113),.res(r90_114),.clk(clk),.wout(w90_114));
	PE pe90_115(.x(x115),.w(w90_114),.acc(r90_114),.res(r90_115),.clk(clk),.wout(w90_115));
	PE pe90_116(.x(x116),.w(w90_115),.acc(r90_115),.res(r90_116),.clk(clk),.wout(w90_116));
	PE pe90_117(.x(x117),.w(w90_116),.acc(r90_116),.res(r90_117),.clk(clk),.wout(w90_117));
	PE pe90_118(.x(x118),.w(w90_117),.acc(r90_117),.res(r90_118),.clk(clk),.wout(w90_118));
	PE pe90_119(.x(x119),.w(w90_118),.acc(r90_118),.res(r90_119),.clk(clk),.wout(w90_119));
	PE pe90_120(.x(x120),.w(w90_119),.acc(r90_119),.res(r90_120),.clk(clk),.wout(w90_120));
	PE pe90_121(.x(x121),.w(w90_120),.acc(r90_120),.res(r90_121),.clk(clk),.wout(w90_121));
	PE pe90_122(.x(x122),.w(w90_121),.acc(r90_121),.res(r90_122),.clk(clk),.wout(w90_122));
	PE pe90_123(.x(x123),.w(w90_122),.acc(r90_122),.res(r90_123),.clk(clk),.wout(w90_123));
	PE pe90_124(.x(x124),.w(w90_123),.acc(r90_123),.res(r90_124),.clk(clk),.wout(w90_124));
	PE pe90_125(.x(x125),.w(w90_124),.acc(r90_124),.res(r90_125),.clk(clk),.wout(w90_125));
	PE pe90_126(.x(x126),.w(w90_125),.acc(r90_125),.res(r90_126),.clk(clk),.wout(w90_126));
	PE pe90_127(.x(x127),.w(w90_126),.acc(r90_126),.res(result90),.clk(clk),.wout(weight90));

	PE pe91_0(.x(x0),.w(w91),.acc(32'h0),.res(r91_0),.clk(clk),.wout(w91_0));
	PE pe91_1(.x(x1),.w(w91_0),.acc(r91_0),.res(r91_1),.clk(clk),.wout(w91_1));
	PE pe91_2(.x(x2),.w(w91_1),.acc(r91_1),.res(r91_2),.clk(clk),.wout(w91_2));
	PE pe91_3(.x(x3),.w(w91_2),.acc(r91_2),.res(r91_3),.clk(clk),.wout(w91_3));
	PE pe91_4(.x(x4),.w(w91_3),.acc(r91_3),.res(r91_4),.clk(clk),.wout(w91_4));
	PE pe91_5(.x(x5),.w(w91_4),.acc(r91_4),.res(r91_5),.clk(clk),.wout(w91_5));
	PE pe91_6(.x(x6),.w(w91_5),.acc(r91_5),.res(r91_6),.clk(clk),.wout(w91_6));
	PE pe91_7(.x(x7),.w(w91_6),.acc(r91_6),.res(r91_7),.clk(clk),.wout(w91_7));
	PE pe91_8(.x(x8),.w(w91_7),.acc(r91_7),.res(r91_8),.clk(clk),.wout(w91_8));
	PE pe91_9(.x(x9),.w(w91_8),.acc(r91_8),.res(r91_9),.clk(clk),.wout(w91_9));
	PE pe91_10(.x(x10),.w(w91_9),.acc(r91_9),.res(r91_10),.clk(clk),.wout(w91_10));
	PE pe91_11(.x(x11),.w(w91_10),.acc(r91_10),.res(r91_11),.clk(clk),.wout(w91_11));
	PE pe91_12(.x(x12),.w(w91_11),.acc(r91_11),.res(r91_12),.clk(clk),.wout(w91_12));
	PE pe91_13(.x(x13),.w(w91_12),.acc(r91_12),.res(r91_13),.clk(clk),.wout(w91_13));
	PE pe91_14(.x(x14),.w(w91_13),.acc(r91_13),.res(r91_14),.clk(clk),.wout(w91_14));
	PE pe91_15(.x(x15),.w(w91_14),.acc(r91_14),.res(r91_15),.clk(clk),.wout(w91_15));
	PE pe91_16(.x(x16),.w(w91_15),.acc(r91_15),.res(r91_16),.clk(clk),.wout(w91_16));
	PE pe91_17(.x(x17),.w(w91_16),.acc(r91_16),.res(r91_17),.clk(clk),.wout(w91_17));
	PE pe91_18(.x(x18),.w(w91_17),.acc(r91_17),.res(r91_18),.clk(clk),.wout(w91_18));
	PE pe91_19(.x(x19),.w(w91_18),.acc(r91_18),.res(r91_19),.clk(clk),.wout(w91_19));
	PE pe91_20(.x(x20),.w(w91_19),.acc(r91_19),.res(r91_20),.clk(clk),.wout(w91_20));
	PE pe91_21(.x(x21),.w(w91_20),.acc(r91_20),.res(r91_21),.clk(clk),.wout(w91_21));
	PE pe91_22(.x(x22),.w(w91_21),.acc(r91_21),.res(r91_22),.clk(clk),.wout(w91_22));
	PE pe91_23(.x(x23),.w(w91_22),.acc(r91_22),.res(r91_23),.clk(clk),.wout(w91_23));
	PE pe91_24(.x(x24),.w(w91_23),.acc(r91_23),.res(r91_24),.clk(clk),.wout(w91_24));
	PE pe91_25(.x(x25),.w(w91_24),.acc(r91_24),.res(r91_25),.clk(clk),.wout(w91_25));
	PE pe91_26(.x(x26),.w(w91_25),.acc(r91_25),.res(r91_26),.clk(clk),.wout(w91_26));
	PE pe91_27(.x(x27),.w(w91_26),.acc(r91_26),.res(r91_27),.clk(clk),.wout(w91_27));
	PE pe91_28(.x(x28),.w(w91_27),.acc(r91_27),.res(r91_28),.clk(clk),.wout(w91_28));
	PE pe91_29(.x(x29),.w(w91_28),.acc(r91_28),.res(r91_29),.clk(clk),.wout(w91_29));
	PE pe91_30(.x(x30),.w(w91_29),.acc(r91_29),.res(r91_30),.clk(clk),.wout(w91_30));
	PE pe91_31(.x(x31),.w(w91_30),.acc(r91_30),.res(r91_31),.clk(clk),.wout(w91_31));
	PE pe91_32(.x(x32),.w(w91_31),.acc(r91_31),.res(r91_32),.clk(clk),.wout(w91_32));
	PE pe91_33(.x(x33),.w(w91_32),.acc(r91_32),.res(r91_33),.clk(clk),.wout(w91_33));
	PE pe91_34(.x(x34),.w(w91_33),.acc(r91_33),.res(r91_34),.clk(clk),.wout(w91_34));
	PE pe91_35(.x(x35),.w(w91_34),.acc(r91_34),.res(r91_35),.clk(clk),.wout(w91_35));
	PE pe91_36(.x(x36),.w(w91_35),.acc(r91_35),.res(r91_36),.clk(clk),.wout(w91_36));
	PE pe91_37(.x(x37),.w(w91_36),.acc(r91_36),.res(r91_37),.clk(clk),.wout(w91_37));
	PE pe91_38(.x(x38),.w(w91_37),.acc(r91_37),.res(r91_38),.clk(clk),.wout(w91_38));
	PE pe91_39(.x(x39),.w(w91_38),.acc(r91_38),.res(r91_39),.clk(clk),.wout(w91_39));
	PE pe91_40(.x(x40),.w(w91_39),.acc(r91_39),.res(r91_40),.clk(clk),.wout(w91_40));
	PE pe91_41(.x(x41),.w(w91_40),.acc(r91_40),.res(r91_41),.clk(clk),.wout(w91_41));
	PE pe91_42(.x(x42),.w(w91_41),.acc(r91_41),.res(r91_42),.clk(clk),.wout(w91_42));
	PE pe91_43(.x(x43),.w(w91_42),.acc(r91_42),.res(r91_43),.clk(clk),.wout(w91_43));
	PE pe91_44(.x(x44),.w(w91_43),.acc(r91_43),.res(r91_44),.clk(clk),.wout(w91_44));
	PE pe91_45(.x(x45),.w(w91_44),.acc(r91_44),.res(r91_45),.clk(clk),.wout(w91_45));
	PE pe91_46(.x(x46),.w(w91_45),.acc(r91_45),.res(r91_46),.clk(clk),.wout(w91_46));
	PE pe91_47(.x(x47),.w(w91_46),.acc(r91_46),.res(r91_47),.clk(clk),.wout(w91_47));
	PE pe91_48(.x(x48),.w(w91_47),.acc(r91_47),.res(r91_48),.clk(clk),.wout(w91_48));
	PE pe91_49(.x(x49),.w(w91_48),.acc(r91_48),.res(r91_49),.clk(clk),.wout(w91_49));
	PE pe91_50(.x(x50),.w(w91_49),.acc(r91_49),.res(r91_50),.clk(clk),.wout(w91_50));
	PE pe91_51(.x(x51),.w(w91_50),.acc(r91_50),.res(r91_51),.clk(clk),.wout(w91_51));
	PE pe91_52(.x(x52),.w(w91_51),.acc(r91_51),.res(r91_52),.clk(clk),.wout(w91_52));
	PE pe91_53(.x(x53),.w(w91_52),.acc(r91_52),.res(r91_53),.clk(clk),.wout(w91_53));
	PE pe91_54(.x(x54),.w(w91_53),.acc(r91_53),.res(r91_54),.clk(clk),.wout(w91_54));
	PE pe91_55(.x(x55),.w(w91_54),.acc(r91_54),.res(r91_55),.clk(clk),.wout(w91_55));
	PE pe91_56(.x(x56),.w(w91_55),.acc(r91_55),.res(r91_56),.clk(clk),.wout(w91_56));
	PE pe91_57(.x(x57),.w(w91_56),.acc(r91_56),.res(r91_57),.clk(clk),.wout(w91_57));
	PE pe91_58(.x(x58),.w(w91_57),.acc(r91_57),.res(r91_58),.clk(clk),.wout(w91_58));
	PE pe91_59(.x(x59),.w(w91_58),.acc(r91_58),.res(r91_59),.clk(clk),.wout(w91_59));
	PE pe91_60(.x(x60),.w(w91_59),.acc(r91_59),.res(r91_60),.clk(clk),.wout(w91_60));
	PE pe91_61(.x(x61),.w(w91_60),.acc(r91_60),.res(r91_61),.clk(clk),.wout(w91_61));
	PE pe91_62(.x(x62),.w(w91_61),.acc(r91_61),.res(r91_62),.clk(clk),.wout(w91_62));
	PE pe91_63(.x(x63),.w(w91_62),.acc(r91_62),.res(r91_63),.clk(clk),.wout(w91_63));
	PE pe91_64(.x(x64),.w(w91_63),.acc(r91_63),.res(r91_64),.clk(clk),.wout(w91_64));
	PE pe91_65(.x(x65),.w(w91_64),.acc(r91_64),.res(r91_65),.clk(clk),.wout(w91_65));
	PE pe91_66(.x(x66),.w(w91_65),.acc(r91_65),.res(r91_66),.clk(clk),.wout(w91_66));
	PE pe91_67(.x(x67),.w(w91_66),.acc(r91_66),.res(r91_67),.clk(clk),.wout(w91_67));
	PE pe91_68(.x(x68),.w(w91_67),.acc(r91_67),.res(r91_68),.clk(clk),.wout(w91_68));
	PE pe91_69(.x(x69),.w(w91_68),.acc(r91_68),.res(r91_69),.clk(clk),.wout(w91_69));
	PE pe91_70(.x(x70),.w(w91_69),.acc(r91_69),.res(r91_70),.clk(clk),.wout(w91_70));
	PE pe91_71(.x(x71),.w(w91_70),.acc(r91_70),.res(r91_71),.clk(clk),.wout(w91_71));
	PE pe91_72(.x(x72),.w(w91_71),.acc(r91_71),.res(r91_72),.clk(clk),.wout(w91_72));
	PE pe91_73(.x(x73),.w(w91_72),.acc(r91_72),.res(r91_73),.clk(clk),.wout(w91_73));
	PE pe91_74(.x(x74),.w(w91_73),.acc(r91_73),.res(r91_74),.clk(clk),.wout(w91_74));
	PE pe91_75(.x(x75),.w(w91_74),.acc(r91_74),.res(r91_75),.clk(clk),.wout(w91_75));
	PE pe91_76(.x(x76),.w(w91_75),.acc(r91_75),.res(r91_76),.clk(clk),.wout(w91_76));
	PE pe91_77(.x(x77),.w(w91_76),.acc(r91_76),.res(r91_77),.clk(clk),.wout(w91_77));
	PE pe91_78(.x(x78),.w(w91_77),.acc(r91_77),.res(r91_78),.clk(clk),.wout(w91_78));
	PE pe91_79(.x(x79),.w(w91_78),.acc(r91_78),.res(r91_79),.clk(clk),.wout(w91_79));
	PE pe91_80(.x(x80),.w(w91_79),.acc(r91_79),.res(r91_80),.clk(clk),.wout(w91_80));
	PE pe91_81(.x(x81),.w(w91_80),.acc(r91_80),.res(r91_81),.clk(clk),.wout(w91_81));
	PE pe91_82(.x(x82),.w(w91_81),.acc(r91_81),.res(r91_82),.clk(clk),.wout(w91_82));
	PE pe91_83(.x(x83),.w(w91_82),.acc(r91_82),.res(r91_83),.clk(clk),.wout(w91_83));
	PE pe91_84(.x(x84),.w(w91_83),.acc(r91_83),.res(r91_84),.clk(clk),.wout(w91_84));
	PE pe91_85(.x(x85),.w(w91_84),.acc(r91_84),.res(r91_85),.clk(clk),.wout(w91_85));
	PE pe91_86(.x(x86),.w(w91_85),.acc(r91_85),.res(r91_86),.clk(clk),.wout(w91_86));
	PE pe91_87(.x(x87),.w(w91_86),.acc(r91_86),.res(r91_87),.clk(clk),.wout(w91_87));
	PE pe91_88(.x(x88),.w(w91_87),.acc(r91_87),.res(r91_88),.clk(clk),.wout(w91_88));
	PE pe91_89(.x(x89),.w(w91_88),.acc(r91_88),.res(r91_89),.clk(clk),.wout(w91_89));
	PE pe91_90(.x(x90),.w(w91_89),.acc(r91_89),.res(r91_90),.clk(clk),.wout(w91_90));
	PE pe91_91(.x(x91),.w(w91_90),.acc(r91_90),.res(r91_91),.clk(clk),.wout(w91_91));
	PE pe91_92(.x(x92),.w(w91_91),.acc(r91_91),.res(r91_92),.clk(clk),.wout(w91_92));
	PE pe91_93(.x(x93),.w(w91_92),.acc(r91_92),.res(r91_93),.clk(clk),.wout(w91_93));
	PE pe91_94(.x(x94),.w(w91_93),.acc(r91_93),.res(r91_94),.clk(clk),.wout(w91_94));
	PE pe91_95(.x(x95),.w(w91_94),.acc(r91_94),.res(r91_95),.clk(clk),.wout(w91_95));
	PE pe91_96(.x(x96),.w(w91_95),.acc(r91_95),.res(r91_96),.clk(clk),.wout(w91_96));
	PE pe91_97(.x(x97),.w(w91_96),.acc(r91_96),.res(r91_97),.clk(clk),.wout(w91_97));
	PE pe91_98(.x(x98),.w(w91_97),.acc(r91_97),.res(r91_98),.clk(clk),.wout(w91_98));
	PE pe91_99(.x(x99),.w(w91_98),.acc(r91_98),.res(r91_99),.clk(clk),.wout(w91_99));
	PE pe91_100(.x(x100),.w(w91_99),.acc(r91_99),.res(r91_100),.clk(clk),.wout(w91_100));
	PE pe91_101(.x(x101),.w(w91_100),.acc(r91_100),.res(r91_101),.clk(clk),.wout(w91_101));
	PE pe91_102(.x(x102),.w(w91_101),.acc(r91_101),.res(r91_102),.clk(clk),.wout(w91_102));
	PE pe91_103(.x(x103),.w(w91_102),.acc(r91_102),.res(r91_103),.clk(clk),.wout(w91_103));
	PE pe91_104(.x(x104),.w(w91_103),.acc(r91_103),.res(r91_104),.clk(clk),.wout(w91_104));
	PE pe91_105(.x(x105),.w(w91_104),.acc(r91_104),.res(r91_105),.clk(clk),.wout(w91_105));
	PE pe91_106(.x(x106),.w(w91_105),.acc(r91_105),.res(r91_106),.clk(clk),.wout(w91_106));
	PE pe91_107(.x(x107),.w(w91_106),.acc(r91_106),.res(r91_107),.clk(clk),.wout(w91_107));
	PE pe91_108(.x(x108),.w(w91_107),.acc(r91_107),.res(r91_108),.clk(clk),.wout(w91_108));
	PE pe91_109(.x(x109),.w(w91_108),.acc(r91_108),.res(r91_109),.clk(clk),.wout(w91_109));
	PE pe91_110(.x(x110),.w(w91_109),.acc(r91_109),.res(r91_110),.clk(clk),.wout(w91_110));
	PE pe91_111(.x(x111),.w(w91_110),.acc(r91_110),.res(r91_111),.clk(clk),.wout(w91_111));
	PE pe91_112(.x(x112),.w(w91_111),.acc(r91_111),.res(r91_112),.clk(clk),.wout(w91_112));
	PE pe91_113(.x(x113),.w(w91_112),.acc(r91_112),.res(r91_113),.clk(clk),.wout(w91_113));
	PE pe91_114(.x(x114),.w(w91_113),.acc(r91_113),.res(r91_114),.clk(clk),.wout(w91_114));
	PE pe91_115(.x(x115),.w(w91_114),.acc(r91_114),.res(r91_115),.clk(clk),.wout(w91_115));
	PE pe91_116(.x(x116),.w(w91_115),.acc(r91_115),.res(r91_116),.clk(clk),.wout(w91_116));
	PE pe91_117(.x(x117),.w(w91_116),.acc(r91_116),.res(r91_117),.clk(clk),.wout(w91_117));
	PE pe91_118(.x(x118),.w(w91_117),.acc(r91_117),.res(r91_118),.clk(clk),.wout(w91_118));
	PE pe91_119(.x(x119),.w(w91_118),.acc(r91_118),.res(r91_119),.clk(clk),.wout(w91_119));
	PE pe91_120(.x(x120),.w(w91_119),.acc(r91_119),.res(r91_120),.clk(clk),.wout(w91_120));
	PE pe91_121(.x(x121),.w(w91_120),.acc(r91_120),.res(r91_121),.clk(clk),.wout(w91_121));
	PE pe91_122(.x(x122),.w(w91_121),.acc(r91_121),.res(r91_122),.clk(clk),.wout(w91_122));
	PE pe91_123(.x(x123),.w(w91_122),.acc(r91_122),.res(r91_123),.clk(clk),.wout(w91_123));
	PE pe91_124(.x(x124),.w(w91_123),.acc(r91_123),.res(r91_124),.clk(clk),.wout(w91_124));
	PE pe91_125(.x(x125),.w(w91_124),.acc(r91_124),.res(r91_125),.clk(clk),.wout(w91_125));
	PE pe91_126(.x(x126),.w(w91_125),.acc(r91_125),.res(r91_126),.clk(clk),.wout(w91_126));
	PE pe91_127(.x(x127),.w(w91_126),.acc(r91_126),.res(result91),.clk(clk),.wout(weight91));

	PE pe92_0(.x(x0),.w(w92),.acc(32'h0),.res(r92_0),.clk(clk),.wout(w92_0));
	PE pe92_1(.x(x1),.w(w92_0),.acc(r92_0),.res(r92_1),.clk(clk),.wout(w92_1));
	PE pe92_2(.x(x2),.w(w92_1),.acc(r92_1),.res(r92_2),.clk(clk),.wout(w92_2));
	PE pe92_3(.x(x3),.w(w92_2),.acc(r92_2),.res(r92_3),.clk(clk),.wout(w92_3));
	PE pe92_4(.x(x4),.w(w92_3),.acc(r92_3),.res(r92_4),.clk(clk),.wout(w92_4));
	PE pe92_5(.x(x5),.w(w92_4),.acc(r92_4),.res(r92_5),.clk(clk),.wout(w92_5));
	PE pe92_6(.x(x6),.w(w92_5),.acc(r92_5),.res(r92_6),.clk(clk),.wout(w92_6));
	PE pe92_7(.x(x7),.w(w92_6),.acc(r92_6),.res(r92_7),.clk(clk),.wout(w92_7));
	PE pe92_8(.x(x8),.w(w92_7),.acc(r92_7),.res(r92_8),.clk(clk),.wout(w92_8));
	PE pe92_9(.x(x9),.w(w92_8),.acc(r92_8),.res(r92_9),.clk(clk),.wout(w92_9));
	PE pe92_10(.x(x10),.w(w92_9),.acc(r92_9),.res(r92_10),.clk(clk),.wout(w92_10));
	PE pe92_11(.x(x11),.w(w92_10),.acc(r92_10),.res(r92_11),.clk(clk),.wout(w92_11));
	PE pe92_12(.x(x12),.w(w92_11),.acc(r92_11),.res(r92_12),.clk(clk),.wout(w92_12));
	PE pe92_13(.x(x13),.w(w92_12),.acc(r92_12),.res(r92_13),.clk(clk),.wout(w92_13));
	PE pe92_14(.x(x14),.w(w92_13),.acc(r92_13),.res(r92_14),.clk(clk),.wout(w92_14));
	PE pe92_15(.x(x15),.w(w92_14),.acc(r92_14),.res(r92_15),.clk(clk),.wout(w92_15));
	PE pe92_16(.x(x16),.w(w92_15),.acc(r92_15),.res(r92_16),.clk(clk),.wout(w92_16));
	PE pe92_17(.x(x17),.w(w92_16),.acc(r92_16),.res(r92_17),.clk(clk),.wout(w92_17));
	PE pe92_18(.x(x18),.w(w92_17),.acc(r92_17),.res(r92_18),.clk(clk),.wout(w92_18));
	PE pe92_19(.x(x19),.w(w92_18),.acc(r92_18),.res(r92_19),.clk(clk),.wout(w92_19));
	PE pe92_20(.x(x20),.w(w92_19),.acc(r92_19),.res(r92_20),.clk(clk),.wout(w92_20));
	PE pe92_21(.x(x21),.w(w92_20),.acc(r92_20),.res(r92_21),.clk(clk),.wout(w92_21));
	PE pe92_22(.x(x22),.w(w92_21),.acc(r92_21),.res(r92_22),.clk(clk),.wout(w92_22));
	PE pe92_23(.x(x23),.w(w92_22),.acc(r92_22),.res(r92_23),.clk(clk),.wout(w92_23));
	PE pe92_24(.x(x24),.w(w92_23),.acc(r92_23),.res(r92_24),.clk(clk),.wout(w92_24));
	PE pe92_25(.x(x25),.w(w92_24),.acc(r92_24),.res(r92_25),.clk(clk),.wout(w92_25));
	PE pe92_26(.x(x26),.w(w92_25),.acc(r92_25),.res(r92_26),.clk(clk),.wout(w92_26));
	PE pe92_27(.x(x27),.w(w92_26),.acc(r92_26),.res(r92_27),.clk(clk),.wout(w92_27));
	PE pe92_28(.x(x28),.w(w92_27),.acc(r92_27),.res(r92_28),.clk(clk),.wout(w92_28));
	PE pe92_29(.x(x29),.w(w92_28),.acc(r92_28),.res(r92_29),.clk(clk),.wout(w92_29));
	PE pe92_30(.x(x30),.w(w92_29),.acc(r92_29),.res(r92_30),.clk(clk),.wout(w92_30));
	PE pe92_31(.x(x31),.w(w92_30),.acc(r92_30),.res(r92_31),.clk(clk),.wout(w92_31));
	PE pe92_32(.x(x32),.w(w92_31),.acc(r92_31),.res(r92_32),.clk(clk),.wout(w92_32));
	PE pe92_33(.x(x33),.w(w92_32),.acc(r92_32),.res(r92_33),.clk(clk),.wout(w92_33));
	PE pe92_34(.x(x34),.w(w92_33),.acc(r92_33),.res(r92_34),.clk(clk),.wout(w92_34));
	PE pe92_35(.x(x35),.w(w92_34),.acc(r92_34),.res(r92_35),.clk(clk),.wout(w92_35));
	PE pe92_36(.x(x36),.w(w92_35),.acc(r92_35),.res(r92_36),.clk(clk),.wout(w92_36));
	PE pe92_37(.x(x37),.w(w92_36),.acc(r92_36),.res(r92_37),.clk(clk),.wout(w92_37));
	PE pe92_38(.x(x38),.w(w92_37),.acc(r92_37),.res(r92_38),.clk(clk),.wout(w92_38));
	PE pe92_39(.x(x39),.w(w92_38),.acc(r92_38),.res(r92_39),.clk(clk),.wout(w92_39));
	PE pe92_40(.x(x40),.w(w92_39),.acc(r92_39),.res(r92_40),.clk(clk),.wout(w92_40));
	PE pe92_41(.x(x41),.w(w92_40),.acc(r92_40),.res(r92_41),.clk(clk),.wout(w92_41));
	PE pe92_42(.x(x42),.w(w92_41),.acc(r92_41),.res(r92_42),.clk(clk),.wout(w92_42));
	PE pe92_43(.x(x43),.w(w92_42),.acc(r92_42),.res(r92_43),.clk(clk),.wout(w92_43));
	PE pe92_44(.x(x44),.w(w92_43),.acc(r92_43),.res(r92_44),.clk(clk),.wout(w92_44));
	PE pe92_45(.x(x45),.w(w92_44),.acc(r92_44),.res(r92_45),.clk(clk),.wout(w92_45));
	PE pe92_46(.x(x46),.w(w92_45),.acc(r92_45),.res(r92_46),.clk(clk),.wout(w92_46));
	PE pe92_47(.x(x47),.w(w92_46),.acc(r92_46),.res(r92_47),.clk(clk),.wout(w92_47));
	PE pe92_48(.x(x48),.w(w92_47),.acc(r92_47),.res(r92_48),.clk(clk),.wout(w92_48));
	PE pe92_49(.x(x49),.w(w92_48),.acc(r92_48),.res(r92_49),.clk(clk),.wout(w92_49));
	PE pe92_50(.x(x50),.w(w92_49),.acc(r92_49),.res(r92_50),.clk(clk),.wout(w92_50));
	PE pe92_51(.x(x51),.w(w92_50),.acc(r92_50),.res(r92_51),.clk(clk),.wout(w92_51));
	PE pe92_52(.x(x52),.w(w92_51),.acc(r92_51),.res(r92_52),.clk(clk),.wout(w92_52));
	PE pe92_53(.x(x53),.w(w92_52),.acc(r92_52),.res(r92_53),.clk(clk),.wout(w92_53));
	PE pe92_54(.x(x54),.w(w92_53),.acc(r92_53),.res(r92_54),.clk(clk),.wout(w92_54));
	PE pe92_55(.x(x55),.w(w92_54),.acc(r92_54),.res(r92_55),.clk(clk),.wout(w92_55));
	PE pe92_56(.x(x56),.w(w92_55),.acc(r92_55),.res(r92_56),.clk(clk),.wout(w92_56));
	PE pe92_57(.x(x57),.w(w92_56),.acc(r92_56),.res(r92_57),.clk(clk),.wout(w92_57));
	PE pe92_58(.x(x58),.w(w92_57),.acc(r92_57),.res(r92_58),.clk(clk),.wout(w92_58));
	PE pe92_59(.x(x59),.w(w92_58),.acc(r92_58),.res(r92_59),.clk(clk),.wout(w92_59));
	PE pe92_60(.x(x60),.w(w92_59),.acc(r92_59),.res(r92_60),.clk(clk),.wout(w92_60));
	PE pe92_61(.x(x61),.w(w92_60),.acc(r92_60),.res(r92_61),.clk(clk),.wout(w92_61));
	PE pe92_62(.x(x62),.w(w92_61),.acc(r92_61),.res(r92_62),.clk(clk),.wout(w92_62));
	PE pe92_63(.x(x63),.w(w92_62),.acc(r92_62),.res(r92_63),.clk(clk),.wout(w92_63));
	PE pe92_64(.x(x64),.w(w92_63),.acc(r92_63),.res(r92_64),.clk(clk),.wout(w92_64));
	PE pe92_65(.x(x65),.w(w92_64),.acc(r92_64),.res(r92_65),.clk(clk),.wout(w92_65));
	PE pe92_66(.x(x66),.w(w92_65),.acc(r92_65),.res(r92_66),.clk(clk),.wout(w92_66));
	PE pe92_67(.x(x67),.w(w92_66),.acc(r92_66),.res(r92_67),.clk(clk),.wout(w92_67));
	PE pe92_68(.x(x68),.w(w92_67),.acc(r92_67),.res(r92_68),.clk(clk),.wout(w92_68));
	PE pe92_69(.x(x69),.w(w92_68),.acc(r92_68),.res(r92_69),.clk(clk),.wout(w92_69));
	PE pe92_70(.x(x70),.w(w92_69),.acc(r92_69),.res(r92_70),.clk(clk),.wout(w92_70));
	PE pe92_71(.x(x71),.w(w92_70),.acc(r92_70),.res(r92_71),.clk(clk),.wout(w92_71));
	PE pe92_72(.x(x72),.w(w92_71),.acc(r92_71),.res(r92_72),.clk(clk),.wout(w92_72));
	PE pe92_73(.x(x73),.w(w92_72),.acc(r92_72),.res(r92_73),.clk(clk),.wout(w92_73));
	PE pe92_74(.x(x74),.w(w92_73),.acc(r92_73),.res(r92_74),.clk(clk),.wout(w92_74));
	PE pe92_75(.x(x75),.w(w92_74),.acc(r92_74),.res(r92_75),.clk(clk),.wout(w92_75));
	PE pe92_76(.x(x76),.w(w92_75),.acc(r92_75),.res(r92_76),.clk(clk),.wout(w92_76));
	PE pe92_77(.x(x77),.w(w92_76),.acc(r92_76),.res(r92_77),.clk(clk),.wout(w92_77));
	PE pe92_78(.x(x78),.w(w92_77),.acc(r92_77),.res(r92_78),.clk(clk),.wout(w92_78));
	PE pe92_79(.x(x79),.w(w92_78),.acc(r92_78),.res(r92_79),.clk(clk),.wout(w92_79));
	PE pe92_80(.x(x80),.w(w92_79),.acc(r92_79),.res(r92_80),.clk(clk),.wout(w92_80));
	PE pe92_81(.x(x81),.w(w92_80),.acc(r92_80),.res(r92_81),.clk(clk),.wout(w92_81));
	PE pe92_82(.x(x82),.w(w92_81),.acc(r92_81),.res(r92_82),.clk(clk),.wout(w92_82));
	PE pe92_83(.x(x83),.w(w92_82),.acc(r92_82),.res(r92_83),.clk(clk),.wout(w92_83));
	PE pe92_84(.x(x84),.w(w92_83),.acc(r92_83),.res(r92_84),.clk(clk),.wout(w92_84));
	PE pe92_85(.x(x85),.w(w92_84),.acc(r92_84),.res(r92_85),.clk(clk),.wout(w92_85));
	PE pe92_86(.x(x86),.w(w92_85),.acc(r92_85),.res(r92_86),.clk(clk),.wout(w92_86));
	PE pe92_87(.x(x87),.w(w92_86),.acc(r92_86),.res(r92_87),.clk(clk),.wout(w92_87));
	PE pe92_88(.x(x88),.w(w92_87),.acc(r92_87),.res(r92_88),.clk(clk),.wout(w92_88));
	PE pe92_89(.x(x89),.w(w92_88),.acc(r92_88),.res(r92_89),.clk(clk),.wout(w92_89));
	PE pe92_90(.x(x90),.w(w92_89),.acc(r92_89),.res(r92_90),.clk(clk),.wout(w92_90));
	PE pe92_91(.x(x91),.w(w92_90),.acc(r92_90),.res(r92_91),.clk(clk),.wout(w92_91));
	PE pe92_92(.x(x92),.w(w92_91),.acc(r92_91),.res(r92_92),.clk(clk),.wout(w92_92));
	PE pe92_93(.x(x93),.w(w92_92),.acc(r92_92),.res(r92_93),.clk(clk),.wout(w92_93));
	PE pe92_94(.x(x94),.w(w92_93),.acc(r92_93),.res(r92_94),.clk(clk),.wout(w92_94));
	PE pe92_95(.x(x95),.w(w92_94),.acc(r92_94),.res(r92_95),.clk(clk),.wout(w92_95));
	PE pe92_96(.x(x96),.w(w92_95),.acc(r92_95),.res(r92_96),.clk(clk),.wout(w92_96));
	PE pe92_97(.x(x97),.w(w92_96),.acc(r92_96),.res(r92_97),.clk(clk),.wout(w92_97));
	PE pe92_98(.x(x98),.w(w92_97),.acc(r92_97),.res(r92_98),.clk(clk),.wout(w92_98));
	PE pe92_99(.x(x99),.w(w92_98),.acc(r92_98),.res(r92_99),.clk(clk),.wout(w92_99));
	PE pe92_100(.x(x100),.w(w92_99),.acc(r92_99),.res(r92_100),.clk(clk),.wout(w92_100));
	PE pe92_101(.x(x101),.w(w92_100),.acc(r92_100),.res(r92_101),.clk(clk),.wout(w92_101));
	PE pe92_102(.x(x102),.w(w92_101),.acc(r92_101),.res(r92_102),.clk(clk),.wout(w92_102));
	PE pe92_103(.x(x103),.w(w92_102),.acc(r92_102),.res(r92_103),.clk(clk),.wout(w92_103));
	PE pe92_104(.x(x104),.w(w92_103),.acc(r92_103),.res(r92_104),.clk(clk),.wout(w92_104));
	PE pe92_105(.x(x105),.w(w92_104),.acc(r92_104),.res(r92_105),.clk(clk),.wout(w92_105));
	PE pe92_106(.x(x106),.w(w92_105),.acc(r92_105),.res(r92_106),.clk(clk),.wout(w92_106));
	PE pe92_107(.x(x107),.w(w92_106),.acc(r92_106),.res(r92_107),.clk(clk),.wout(w92_107));
	PE pe92_108(.x(x108),.w(w92_107),.acc(r92_107),.res(r92_108),.clk(clk),.wout(w92_108));
	PE pe92_109(.x(x109),.w(w92_108),.acc(r92_108),.res(r92_109),.clk(clk),.wout(w92_109));
	PE pe92_110(.x(x110),.w(w92_109),.acc(r92_109),.res(r92_110),.clk(clk),.wout(w92_110));
	PE pe92_111(.x(x111),.w(w92_110),.acc(r92_110),.res(r92_111),.clk(clk),.wout(w92_111));
	PE pe92_112(.x(x112),.w(w92_111),.acc(r92_111),.res(r92_112),.clk(clk),.wout(w92_112));
	PE pe92_113(.x(x113),.w(w92_112),.acc(r92_112),.res(r92_113),.clk(clk),.wout(w92_113));
	PE pe92_114(.x(x114),.w(w92_113),.acc(r92_113),.res(r92_114),.clk(clk),.wout(w92_114));
	PE pe92_115(.x(x115),.w(w92_114),.acc(r92_114),.res(r92_115),.clk(clk),.wout(w92_115));
	PE pe92_116(.x(x116),.w(w92_115),.acc(r92_115),.res(r92_116),.clk(clk),.wout(w92_116));
	PE pe92_117(.x(x117),.w(w92_116),.acc(r92_116),.res(r92_117),.clk(clk),.wout(w92_117));
	PE pe92_118(.x(x118),.w(w92_117),.acc(r92_117),.res(r92_118),.clk(clk),.wout(w92_118));
	PE pe92_119(.x(x119),.w(w92_118),.acc(r92_118),.res(r92_119),.clk(clk),.wout(w92_119));
	PE pe92_120(.x(x120),.w(w92_119),.acc(r92_119),.res(r92_120),.clk(clk),.wout(w92_120));
	PE pe92_121(.x(x121),.w(w92_120),.acc(r92_120),.res(r92_121),.clk(clk),.wout(w92_121));
	PE pe92_122(.x(x122),.w(w92_121),.acc(r92_121),.res(r92_122),.clk(clk),.wout(w92_122));
	PE pe92_123(.x(x123),.w(w92_122),.acc(r92_122),.res(r92_123),.clk(clk),.wout(w92_123));
	PE pe92_124(.x(x124),.w(w92_123),.acc(r92_123),.res(r92_124),.clk(clk),.wout(w92_124));
	PE pe92_125(.x(x125),.w(w92_124),.acc(r92_124),.res(r92_125),.clk(clk),.wout(w92_125));
	PE pe92_126(.x(x126),.w(w92_125),.acc(r92_125),.res(r92_126),.clk(clk),.wout(w92_126));
	PE pe92_127(.x(x127),.w(w92_126),.acc(r92_126),.res(result92),.clk(clk),.wout(weight92));

	PE pe93_0(.x(x0),.w(w93),.acc(32'h0),.res(r93_0),.clk(clk),.wout(w93_0));
	PE pe93_1(.x(x1),.w(w93_0),.acc(r93_0),.res(r93_1),.clk(clk),.wout(w93_1));
	PE pe93_2(.x(x2),.w(w93_1),.acc(r93_1),.res(r93_2),.clk(clk),.wout(w93_2));
	PE pe93_3(.x(x3),.w(w93_2),.acc(r93_2),.res(r93_3),.clk(clk),.wout(w93_3));
	PE pe93_4(.x(x4),.w(w93_3),.acc(r93_3),.res(r93_4),.clk(clk),.wout(w93_4));
	PE pe93_5(.x(x5),.w(w93_4),.acc(r93_4),.res(r93_5),.clk(clk),.wout(w93_5));
	PE pe93_6(.x(x6),.w(w93_5),.acc(r93_5),.res(r93_6),.clk(clk),.wout(w93_6));
	PE pe93_7(.x(x7),.w(w93_6),.acc(r93_6),.res(r93_7),.clk(clk),.wout(w93_7));
	PE pe93_8(.x(x8),.w(w93_7),.acc(r93_7),.res(r93_8),.clk(clk),.wout(w93_8));
	PE pe93_9(.x(x9),.w(w93_8),.acc(r93_8),.res(r93_9),.clk(clk),.wout(w93_9));
	PE pe93_10(.x(x10),.w(w93_9),.acc(r93_9),.res(r93_10),.clk(clk),.wout(w93_10));
	PE pe93_11(.x(x11),.w(w93_10),.acc(r93_10),.res(r93_11),.clk(clk),.wout(w93_11));
	PE pe93_12(.x(x12),.w(w93_11),.acc(r93_11),.res(r93_12),.clk(clk),.wout(w93_12));
	PE pe93_13(.x(x13),.w(w93_12),.acc(r93_12),.res(r93_13),.clk(clk),.wout(w93_13));
	PE pe93_14(.x(x14),.w(w93_13),.acc(r93_13),.res(r93_14),.clk(clk),.wout(w93_14));
	PE pe93_15(.x(x15),.w(w93_14),.acc(r93_14),.res(r93_15),.clk(clk),.wout(w93_15));
	PE pe93_16(.x(x16),.w(w93_15),.acc(r93_15),.res(r93_16),.clk(clk),.wout(w93_16));
	PE pe93_17(.x(x17),.w(w93_16),.acc(r93_16),.res(r93_17),.clk(clk),.wout(w93_17));
	PE pe93_18(.x(x18),.w(w93_17),.acc(r93_17),.res(r93_18),.clk(clk),.wout(w93_18));
	PE pe93_19(.x(x19),.w(w93_18),.acc(r93_18),.res(r93_19),.clk(clk),.wout(w93_19));
	PE pe93_20(.x(x20),.w(w93_19),.acc(r93_19),.res(r93_20),.clk(clk),.wout(w93_20));
	PE pe93_21(.x(x21),.w(w93_20),.acc(r93_20),.res(r93_21),.clk(clk),.wout(w93_21));
	PE pe93_22(.x(x22),.w(w93_21),.acc(r93_21),.res(r93_22),.clk(clk),.wout(w93_22));
	PE pe93_23(.x(x23),.w(w93_22),.acc(r93_22),.res(r93_23),.clk(clk),.wout(w93_23));
	PE pe93_24(.x(x24),.w(w93_23),.acc(r93_23),.res(r93_24),.clk(clk),.wout(w93_24));
	PE pe93_25(.x(x25),.w(w93_24),.acc(r93_24),.res(r93_25),.clk(clk),.wout(w93_25));
	PE pe93_26(.x(x26),.w(w93_25),.acc(r93_25),.res(r93_26),.clk(clk),.wout(w93_26));
	PE pe93_27(.x(x27),.w(w93_26),.acc(r93_26),.res(r93_27),.clk(clk),.wout(w93_27));
	PE pe93_28(.x(x28),.w(w93_27),.acc(r93_27),.res(r93_28),.clk(clk),.wout(w93_28));
	PE pe93_29(.x(x29),.w(w93_28),.acc(r93_28),.res(r93_29),.clk(clk),.wout(w93_29));
	PE pe93_30(.x(x30),.w(w93_29),.acc(r93_29),.res(r93_30),.clk(clk),.wout(w93_30));
	PE pe93_31(.x(x31),.w(w93_30),.acc(r93_30),.res(r93_31),.clk(clk),.wout(w93_31));
	PE pe93_32(.x(x32),.w(w93_31),.acc(r93_31),.res(r93_32),.clk(clk),.wout(w93_32));
	PE pe93_33(.x(x33),.w(w93_32),.acc(r93_32),.res(r93_33),.clk(clk),.wout(w93_33));
	PE pe93_34(.x(x34),.w(w93_33),.acc(r93_33),.res(r93_34),.clk(clk),.wout(w93_34));
	PE pe93_35(.x(x35),.w(w93_34),.acc(r93_34),.res(r93_35),.clk(clk),.wout(w93_35));
	PE pe93_36(.x(x36),.w(w93_35),.acc(r93_35),.res(r93_36),.clk(clk),.wout(w93_36));
	PE pe93_37(.x(x37),.w(w93_36),.acc(r93_36),.res(r93_37),.clk(clk),.wout(w93_37));
	PE pe93_38(.x(x38),.w(w93_37),.acc(r93_37),.res(r93_38),.clk(clk),.wout(w93_38));
	PE pe93_39(.x(x39),.w(w93_38),.acc(r93_38),.res(r93_39),.clk(clk),.wout(w93_39));
	PE pe93_40(.x(x40),.w(w93_39),.acc(r93_39),.res(r93_40),.clk(clk),.wout(w93_40));
	PE pe93_41(.x(x41),.w(w93_40),.acc(r93_40),.res(r93_41),.clk(clk),.wout(w93_41));
	PE pe93_42(.x(x42),.w(w93_41),.acc(r93_41),.res(r93_42),.clk(clk),.wout(w93_42));
	PE pe93_43(.x(x43),.w(w93_42),.acc(r93_42),.res(r93_43),.clk(clk),.wout(w93_43));
	PE pe93_44(.x(x44),.w(w93_43),.acc(r93_43),.res(r93_44),.clk(clk),.wout(w93_44));
	PE pe93_45(.x(x45),.w(w93_44),.acc(r93_44),.res(r93_45),.clk(clk),.wout(w93_45));
	PE pe93_46(.x(x46),.w(w93_45),.acc(r93_45),.res(r93_46),.clk(clk),.wout(w93_46));
	PE pe93_47(.x(x47),.w(w93_46),.acc(r93_46),.res(r93_47),.clk(clk),.wout(w93_47));
	PE pe93_48(.x(x48),.w(w93_47),.acc(r93_47),.res(r93_48),.clk(clk),.wout(w93_48));
	PE pe93_49(.x(x49),.w(w93_48),.acc(r93_48),.res(r93_49),.clk(clk),.wout(w93_49));
	PE pe93_50(.x(x50),.w(w93_49),.acc(r93_49),.res(r93_50),.clk(clk),.wout(w93_50));
	PE pe93_51(.x(x51),.w(w93_50),.acc(r93_50),.res(r93_51),.clk(clk),.wout(w93_51));
	PE pe93_52(.x(x52),.w(w93_51),.acc(r93_51),.res(r93_52),.clk(clk),.wout(w93_52));
	PE pe93_53(.x(x53),.w(w93_52),.acc(r93_52),.res(r93_53),.clk(clk),.wout(w93_53));
	PE pe93_54(.x(x54),.w(w93_53),.acc(r93_53),.res(r93_54),.clk(clk),.wout(w93_54));
	PE pe93_55(.x(x55),.w(w93_54),.acc(r93_54),.res(r93_55),.clk(clk),.wout(w93_55));
	PE pe93_56(.x(x56),.w(w93_55),.acc(r93_55),.res(r93_56),.clk(clk),.wout(w93_56));
	PE pe93_57(.x(x57),.w(w93_56),.acc(r93_56),.res(r93_57),.clk(clk),.wout(w93_57));
	PE pe93_58(.x(x58),.w(w93_57),.acc(r93_57),.res(r93_58),.clk(clk),.wout(w93_58));
	PE pe93_59(.x(x59),.w(w93_58),.acc(r93_58),.res(r93_59),.clk(clk),.wout(w93_59));
	PE pe93_60(.x(x60),.w(w93_59),.acc(r93_59),.res(r93_60),.clk(clk),.wout(w93_60));
	PE pe93_61(.x(x61),.w(w93_60),.acc(r93_60),.res(r93_61),.clk(clk),.wout(w93_61));
	PE pe93_62(.x(x62),.w(w93_61),.acc(r93_61),.res(r93_62),.clk(clk),.wout(w93_62));
	PE pe93_63(.x(x63),.w(w93_62),.acc(r93_62),.res(r93_63),.clk(clk),.wout(w93_63));
	PE pe93_64(.x(x64),.w(w93_63),.acc(r93_63),.res(r93_64),.clk(clk),.wout(w93_64));
	PE pe93_65(.x(x65),.w(w93_64),.acc(r93_64),.res(r93_65),.clk(clk),.wout(w93_65));
	PE pe93_66(.x(x66),.w(w93_65),.acc(r93_65),.res(r93_66),.clk(clk),.wout(w93_66));
	PE pe93_67(.x(x67),.w(w93_66),.acc(r93_66),.res(r93_67),.clk(clk),.wout(w93_67));
	PE pe93_68(.x(x68),.w(w93_67),.acc(r93_67),.res(r93_68),.clk(clk),.wout(w93_68));
	PE pe93_69(.x(x69),.w(w93_68),.acc(r93_68),.res(r93_69),.clk(clk),.wout(w93_69));
	PE pe93_70(.x(x70),.w(w93_69),.acc(r93_69),.res(r93_70),.clk(clk),.wout(w93_70));
	PE pe93_71(.x(x71),.w(w93_70),.acc(r93_70),.res(r93_71),.clk(clk),.wout(w93_71));
	PE pe93_72(.x(x72),.w(w93_71),.acc(r93_71),.res(r93_72),.clk(clk),.wout(w93_72));
	PE pe93_73(.x(x73),.w(w93_72),.acc(r93_72),.res(r93_73),.clk(clk),.wout(w93_73));
	PE pe93_74(.x(x74),.w(w93_73),.acc(r93_73),.res(r93_74),.clk(clk),.wout(w93_74));
	PE pe93_75(.x(x75),.w(w93_74),.acc(r93_74),.res(r93_75),.clk(clk),.wout(w93_75));
	PE pe93_76(.x(x76),.w(w93_75),.acc(r93_75),.res(r93_76),.clk(clk),.wout(w93_76));
	PE pe93_77(.x(x77),.w(w93_76),.acc(r93_76),.res(r93_77),.clk(clk),.wout(w93_77));
	PE pe93_78(.x(x78),.w(w93_77),.acc(r93_77),.res(r93_78),.clk(clk),.wout(w93_78));
	PE pe93_79(.x(x79),.w(w93_78),.acc(r93_78),.res(r93_79),.clk(clk),.wout(w93_79));
	PE pe93_80(.x(x80),.w(w93_79),.acc(r93_79),.res(r93_80),.clk(clk),.wout(w93_80));
	PE pe93_81(.x(x81),.w(w93_80),.acc(r93_80),.res(r93_81),.clk(clk),.wout(w93_81));
	PE pe93_82(.x(x82),.w(w93_81),.acc(r93_81),.res(r93_82),.clk(clk),.wout(w93_82));
	PE pe93_83(.x(x83),.w(w93_82),.acc(r93_82),.res(r93_83),.clk(clk),.wout(w93_83));
	PE pe93_84(.x(x84),.w(w93_83),.acc(r93_83),.res(r93_84),.clk(clk),.wout(w93_84));
	PE pe93_85(.x(x85),.w(w93_84),.acc(r93_84),.res(r93_85),.clk(clk),.wout(w93_85));
	PE pe93_86(.x(x86),.w(w93_85),.acc(r93_85),.res(r93_86),.clk(clk),.wout(w93_86));
	PE pe93_87(.x(x87),.w(w93_86),.acc(r93_86),.res(r93_87),.clk(clk),.wout(w93_87));
	PE pe93_88(.x(x88),.w(w93_87),.acc(r93_87),.res(r93_88),.clk(clk),.wout(w93_88));
	PE pe93_89(.x(x89),.w(w93_88),.acc(r93_88),.res(r93_89),.clk(clk),.wout(w93_89));
	PE pe93_90(.x(x90),.w(w93_89),.acc(r93_89),.res(r93_90),.clk(clk),.wout(w93_90));
	PE pe93_91(.x(x91),.w(w93_90),.acc(r93_90),.res(r93_91),.clk(clk),.wout(w93_91));
	PE pe93_92(.x(x92),.w(w93_91),.acc(r93_91),.res(r93_92),.clk(clk),.wout(w93_92));
	PE pe93_93(.x(x93),.w(w93_92),.acc(r93_92),.res(r93_93),.clk(clk),.wout(w93_93));
	PE pe93_94(.x(x94),.w(w93_93),.acc(r93_93),.res(r93_94),.clk(clk),.wout(w93_94));
	PE pe93_95(.x(x95),.w(w93_94),.acc(r93_94),.res(r93_95),.clk(clk),.wout(w93_95));
	PE pe93_96(.x(x96),.w(w93_95),.acc(r93_95),.res(r93_96),.clk(clk),.wout(w93_96));
	PE pe93_97(.x(x97),.w(w93_96),.acc(r93_96),.res(r93_97),.clk(clk),.wout(w93_97));
	PE pe93_98(.x(x98),.w(w93_97),.acc(r93_97),.res(r93_98),.clk(clk),.wout(w93_98));
	PE pe93_99(.x(x99),.w(w93_98),.acc(r93_98),.res(r93_99),.clk(clk),.wout(w93_99));
	PE pe93_100(.x(x100),.w(w93_99),.acc(r93_99),.res(r93_100),.clk(clk),.wout(w93_100));
	PE pe93_101(.x(x101),.w(w93_100),.acc(r93_100),.res(r93_101),.clk(clk),.wout(w93_101));
	PE pe93_102(.x(x102),.w(w93_101),.acc(r93_101),.res(r93_102),.clk(clk),.wout(w93_102));
	PE pe93_103(.x(x103),.w(w93_102),.acc(r93_102),.res(r93_103),.clk(clk),.wout(w93_103));
	PE pe93_104(.x(x104),.w(w93_103),.acc(r93_103),.res(r93_104),.clk(clk),.wout(w93_104));
	PE pe93_105(.x(x105),.w(w93_104),.acc(r93_104),.res(r93_105),.clk(clk),.wout(w93_105));
	PE pe93_106(.x(x106),.w(w93_105),.acc(r93_105),.res(r93_106),.clk(clk),.wout(w93_106));
	PE pe93_107(.x(x107),.w(w93_106),.acc(r93_106),.res(r93_107),.clk(clk),.wout(w93_107));
	PE pe93_108(.x(x108),.w(w93_107),.acc(r93_107),.res(r93_108),.clk(clk),.wout(w93_108));
	PE pe93_109(.x(x109),.w(w93_108),.acc(r93_108),.res(r93_109),.clk(clk),.wout(w93_109));
	PE pe93_110(.x(x110),.w(w93_109),.acc(r93_109),.res(r93_110),.clk(clk),.wout(w93_110));
	PE pe93_111(.x(x111),.w(w93_110),.acc(r93_110),.res(r93_111),.clk(clk),.wout(w93_111));
	PE pe93_112(.x(x112),.w(w93_111),.acc(r93_111),.res(r93_112),.clk(clk),.wout(w93_112));
	PE pe93_113(.x(x113),.w(w93_112),.acc(r93_112),.res(r93_113),.clk(clk),.wout(w93_113));
	PE pe93_114(.x(x114),.w(w93_113),.acc(r93_113),.res(r93_114),.clk(clk),.wout(w93_114));
	PE pe93_115(.x(x115),.w(w93_114),.acc(r93_114),.res(r93_115),.clk(clk),.wout(w93_115));
	PE pe93_116(.x(x116),.w(w93_115),.acc(r93_115),.res(r93_116),.clk(clk),.wout(w93_116));
	PE pe93_117(.x(x117),.w(w93_116),.acc(r93_116),.res(r93_117),.clk(clk),.wout(w93_117));
	PE pe93_118(.x(x118),.w(w93_117),.acc(r93_117),.res(r93_118),.clk(clk),.wout(w93_118));
	PE pe93_119(.x(x119),.w(w93_118),.acc(r93_118),.res(r93_119),.clk(clk),.wout(w93_119));
	PE pe93_120(.x(x120),.w(w93_119),.acc(r93_119),.res(r93_120),.clk(clk),.wout(w93_120));
	PE pe93_121(.x(x121),.w(w93_120),.acc(r93_120),.res(r93_121),.clk(clk),.wout(w93_121));
	PE pe93_122(.x(x122),.w(w93_121),.acc(r93_121),.res(r93_122),.clk(clk),.wout(w93_122));
	PE pe93_123(.x(x123),.w(w93_122),.acc(r93_122),.res(r93_123),.clk(clk),.wout(w93_123));
	PE pe93_124(.x(x124),.w(w93_123),.acc(r93_123),.res(r93_124),.clk(clk),.wout(w93_124));
	PE pe93_125(.x(x125),.w(w93_124),.acc(r93_124),.res(r93_125),.clk(clk),.wout(w93_125));
	PE pe93_126(.x(x126),.w(w93_125),.acc(r93_125),.res(r93_126),.clk(clk),.wout(w93_126));
	PE pe93_127(.x(x127),.w(w93_126),.acc(r93_126),.res(result93),.clk(clk),.wout(weight93));

	PE pe94_0(.x(x0),.w(w94),.acc(32'h0),.res(r94_0),.clk(clk),.wout(w94_0));
	PE pe94_1(.x(x1),.w(w94_0),.acc(r94_0),.res(r94_1),.clk(clk),.wout(w94_1));
	PE pe94_2(.x(x2),.w(w94_1),.acc(r94_1),.res(r94_2),.clk(clk),.wout(w94_2));
	PE pe94_3(.x(x3),.w(w94_2),.acc(r94_2),.res(r94_3),.clk(clk),.wout(w94_3));
	PE pe94_4(.x(x4),.w(w94_3),.acc(r94_3),.res(r94_4),.clk(clk),.wout(w94_4));
	PE pe94_5(.x(x5),.w(w94_4),.acc(r94_4),.res(r94_5),.clk(clk),.wout(w94_5));
	PE pe94_6(.x(x6),.w(w94_5),.acc(r94_5),.res(r94_6),.clk(clk),.wout(w94_6));
	PE pe94_7(.x(x7),.w(w94_6),.acc(r94_6),.res(r94_7),.clk(clk),.wout(w94_7));
	PE pe94_8(.x(x8),.w(w94_7),.acc(r94_7),.res(r94_8),.clk(clk),.wout(w94_8));
	PE pe94_9(.x(x9),.w(w94_8),.acc(r94_8),.res(r94_9),.clk(clk),.wout(w94_9));
	PE pe94_10(.x(x10),.w(w94_9),.acc(r94_9),.res(r94_10),.clk(clk),.wout(w94_10));
	PE pe94_11(.x(x11),.w(w94_10),.acc(r94_10),.res(r94_11),.clk(clk),.wout(w94_11));
	PE pe94_12(.x(x12),.w(w94_11),.acc(r94_11),.res(r94_12),.clk(clk),.wout(w94_12));
	PE pe94_13(.x(x13),.w(w94_12),.acc(r94_12),.res(r94_13),.clk(clk),.wout(w94_13));
	PE pe94_14(.x(x14),.w(w94_13),.acc(r94_13),.res(r94_14),.clk(clk),.wout(w94_14));
	PE pe94_15(.x(x15),.w(w94_14),.acc(r94_14),.res(r94_15),.clk(clk),.wout(w94_15));
	PE pe94_16(.x(x16),.w(w94_15),.acc(r94_15),.res(r94_16),.clk(clk),.wout(w94_16));
	PE pe94_17(.x(x17),.w(w94_16),.acc(r94_16),.res(r94_17),.clk(clk),.wout(w94_17));
	PE pe94_18(.x(x18),.w(w94_17),.acc(r94_17),.res(r94_18),.clk(clk),.wout(w94_18));
	PE pe94_19(.x(x19),.w(w94_18),.acc(r94_18),.res(r94_19),.clk(clk),.wout(w94_19));
	PE pe94_20(.x(x20),.w(w94_19),.acc(r94_19),.res(r94_20),.clk(clk),.wout(w94_20));
	PE pe94_21(.x(x21),.w(w94_20),.acc(r94_20),.res(r94_21),.clk(clk),.wout(w94_21));
	PE pe94_22(.x(x22),.w(w94_21),.acc(r94_21),.res(r94_22),.clk(clk),.wout(w94_22));
	PE pe94_23(.x(x23),.w(w94_22),.acc(r94_22),.res(r94_23),.clk(clk),.wout(w94_23));
	PE pe94_24(.x(x24),.w(w94_23),.acc(r94_23),.res(r94_24),.clk(clk),.wout(w94_24));
	PE pe94_25(.x(x25),.w(w94_24),.acc(r94_24),.res(r94_25),.clk(clk),.wout(w94_25));
	PE pe94_26(.x(x26),.w(w94_25),.acc(r94_25),.res(r94_26),.clk(clk),.wout(w94_26));
	PE pe94_27(.x(x27),.w(w94_26),.acc(r94_26),.res(r94_27),.clk(clk),.wout(w94_27));
	PE pe94_28(.x(x28),.w(w94_27),.acc(r94_27),.res(r94_28),.clk(clk),.wout(w94_28));
	PE pe94_29(.x(x29),.w(w94_28),.acc(r94_28),.res(r94_29),.clk(clk),.wout(w94_29));
	PE pe94_30(.x(x30),.w(w94_29),.acc(r94_29),.res(r94_30),.clk(clk),.wout(w94_30));
	PE pe94_31(.x(x31),.w(w94_30),.acc(r94_30),.res(r94_31),.clk(clk),.wout(w94_31));
	PE pe94_32(.x(x32),.w(w94_31),.acc(r94_31),.res(r94_32),.clk(clk),.wout(w94_32));
	PE pe94_33(.x(x33),.w(w94_32),.acc(r94_32),.res(r94_33),.clk(clk),.wout(w94_33));
	PE pe94_34(.x(x34),.w(w94_33),.acc(r94_33),.res(r94_34),.clk(clk),.wout(w94_34));
	PE pe94_35(.x(x35),.w(w94_34),.acc(r94_34),.res(r94_35),.clk(clk),.wout(w94_35));
	PE pe94_36(.x(x36),.w(w94_35),.acc(r94_35),.res(r94_36),.clk(clk),.wout(w94_36));
	PE pe94_37(.x(x37),.w(w94_36),.acc(r94_36),.res(r94_37),.clk(clk),.wout(w94_37));
	PE pe94_38(.x(x38),.w(w94_37),.acc(r94_37),.res(r94_38),.clk(clk),.wout(w94_38));
	PE pe94_39(.x(x39),.w(w94_38),.acc(r94_38),.res(r94_39),.clk(clk),.wout(w94_39));
	PE pe94_40(.x(x40),.w(w94_39),.acc(r94_39),.res(r94_40),.clk(clk),.wout(w94_40));
	PE pe94_41(.x(x41),.w(w94_40),.acc(r94_40),.res(r94_41),.clk(clk),.wout(w94_41));
	PE pe94_42(.x(x42),.w(w94_41),.acc(r94_41),.res(r94_42),.clk(clk),.wout(w94_42));
	PE pe94_43(.x(x43),.w(w94_42),.acc(r94_42),.res(r94_43),.clk(clk),.wout(w94_43));
	PE pe94_44(.x(x44),.w(w94_43),.acc(r94_43),.res(r94_44),.clk(clk),.wout(w94_44));
	PE pe94_45(.x(x45),.w(w94_44),.acc(r94_44),.res(r94_45),.clk(clk),.wout(w94_45));
	PE pe94_46(.x(x46),.w(w94_45),.acc(r94_45),.res(r94_46),.clk(clk),.wout(w94_46));
	PE pe94_47(.x(x47),.w(w94_46),.acc(r94_46),.res(r94_47),.clk(clk),.wout(w94_47));
	PE pe94_48(.x(x48),.w(w94_47),.acc(r94_47),.res(r94_48),.clk(clk),.wout(w94_48));
	PE pe94_49(.x(x49),.w(w94_48),.acc(r94_48),.res(r94_49),.clk(clk),.wout(w94_49));
	PE pe94_50(.x(x50),.w(w94_49),.acc(r94_49),.res(r94_50),.clk(clk),.wout(w94_50));
	PE pe94_51(.x(x51),.w(w94_50),.acc(r94_50),.res(r94_51),.clk(clk),.wout(w94_51));
	PE pe94_52(.x(x52),.w(w94_51),.acc(r94_51),.res(r94_52),.clk(clk),.wout(w94_52));
	PE pe94_53(.x(x53),.w(w94_52),.acc(r94_52),.res(r94_53),.clk(clk),.wout(w94_53));
	PE pe94_54(.x(x54),.w(w94_53),.acc(r94_53),.res(r94_54),.clk(clk),.wout(w94_54));
	PE pe94_55(.x(x55),.w(w94_54),.acc(r94_54),.res(r94_55),.clk(clk),.wout(w94_55));
	PE pe94_56(.x(x56),.w(w94_55),.acc(r94_55),.res(r94_56),.clk(clk),.wout(w94_56));
	PE pe94_57(.x(x57),.w(w94_56),.acc(r94_56),.res(r94_57),.clk(clk),.wout(w94_57));
	PE pe94_58(.x(x58),.w(w94_57),.acc(r94_57),.res(r94_58),.clk(clk),.wout(w94_58));
	PE pe94_59(.x(x59),.w(w94_58),.acc(r94_58),.res(r94_59),.clk(clk),.wout(w94_59));
	PE pe94_60(.x(x60),.w(w94_59),.acc(r94_59),.res(r94_60),.clk(clk),.wout(w94_60));
	PE pe94_61(.x(x61),.w(w94_60),.acc(r94_60),.res(r94_61),.clk(clk),.wout(w94_61));
	PE pe94_62(.x(x62),.w(w94_61),.acc(r94_61),.res(r94_62),.clk(clk),.wout(w94_62));
	PE pe94_63(.x(x63),.w(w94_62),.acc(r94_62),.res(r94_63),.clk(clk),.wout(w94_63));
	PE pe94_64(.x(x64),.w(w94_63),.acc(r94_63),.res(r94_64),.clk(clk),.wout(w94_64));
	PE pe94_65(.x(x65),.w(w94_64),.acc(r94_64),.res(r94_65),.clk(clk),.wout(w94_65));
	PE pe94_66(.x(x66),.w(w94_65),.acc(r94_65),.res(r94_66),.clk(clk),.wout(w94_66));
	PE pe94_67(.x(x67),.w(w94_66),.acc(r94_66),.res(r94_67),.clk(clk),.wout(w94_67));
	PE pe94_68(.x(x68),.w(w94_67),.acc(r94_67),.res(r94_68),.clk(clk),.wout(w94_68));
	PE pe94_69(.x(x69),.w(w94_68),.acc(r94_68),.res(r94_69),.clk(clk),.wout(w94_69));
	PE pe94_70(.x(x70),.w(w94_69),.acc(r94_69),.res(r94_70),.clk(clk),.wout(w94_70));
	PE pe94_71(.x(x71),.w(w94_70),.acc(r94_70),.res(r94_71),.clk(clk),.wout(w94_71));
	PE pe94_72(.x(x72),.w(w94_71),.acc(r94_71),.res(r94_72),.clk(clk),.wout(w94_72));
	PE pe94_73(.x(x73),.w(w94_72),.acc(r94_72),.res(r94_73),.clk(clk),.wout(w94_73));
	PE pe94_74(.x(x74),.w(w94_73),.acc(r94_73),.res(r94_74),.clk(clk),.wout(w94_74));
	PE pe94_75(.x(x75),.w(w94_74),.acc(r94_74),.res(r94_75),.clk(clk),.wout(w94_75));
	PE pe94_76(.x(x76),.w(w94_75),.acc(r94_75),.res(r94_76),.clk(clk),.wout(w94_76));
	PE pe94_77(.x(x77),.w(w94_76),.acc(r94_76),.res(r94_77),.clk(clk),.wout(w94_77));
	PE pe94_78(.x(x78),.w(w94_77),.acc(r94_77),.res(r94_78),.clk(clk),.wout(w94_78));
	PE pe94_79(.x(x79),.w(w94_78),.acc(r94_78),.res(r94_79),.clk(clk),.wout(w94_79));
	PE pe94_80(.x(x80),.w(w94_79),.acc(r94_79),.res(r94_80),.clk(clk),.wout(w94_80));
	PE pe94_81(.x(x81),.w(w94_80),.acc(r94_80),.res(r94_81),.clk(clk),.wout(w94_81));
	PE pe94_82(.x(x82),.w(w94_81),.acc(r94_81),.res(r94_82),.clk(clk),.wout(w94_82));
	PE pe94_83(.x(x83),.w(w94_82),.acc(r94_82),.res(r94_83),.clk(clk),.wout(w94_83));
	PE pe94_84(.x(x84),.w(w94_83),.acc(r94_83),.res(r94_84),.clk(clk),.wout(w94_84));
	PE pe94_85(.x(x85),.w(w94_84),.acc(r94_84),.res(r94_85),.clk(clk),.wout(w94_85));
	PE pe94_86(.x(x86),.w(w94_85),.acc(r94_85),.res(r94_86),.clk(clk),.wout(w94_86));
	PE pe94_87(.x(x87),.w(w94_86),.acc(r94_86),.res(r94_87),.clk(clk),.wout(w94_87));
	PE pe94_88(.x(x88),.w(w94_87),.acc(r94_87),.res(r94_88),.clk(clk),.wout(w94_88));
	PE pe94_89(.x(x89),.w(w94_88),.acc(r94_88),.res(r94_89),.clk(clk),.wout(w94_89));
	PE pe94_90(.x(x90),.w(w94_89),.acc(r94_89),.res(r94_90),.clk(clk),.wout(w94_90));
	PE pe94_91(.x(x91),.w(w94_90),.acc(r94_90),.res(r94_91),.clk(clk),.wout(w94_91));
	PE pe94_92(.x(x92),.w(w94_91),.acc(r94_91),.res(r94_92),.clk(clk),.wout(w94_92));
	PE pe94_93(.x(x93),.w(w94_92),.acc(r94_92),.res(r94_93),.clk(clk),.wout(w94_93));
	PE pe94_94(.x(x94),.w(w94_93),.acc(r94_93),.res(r94_94),.clk(clk),.wout(w94_94));
	PE pe94_95(.x(x95),.w(w94_94),.acc(r94_94),.res(r94_95),.clk(clk),.wout(w94_95));
	PE pe94_96(.x(x96),.w(w94_95),.acc(r94_95),.res(r94_96),.clk(clk),.wout(w94_96));
	PE pe94_97(.x(x97),.w(w94_96),.acc(r94_96),.res(r94_97),.clk(clk),.wout(w94_97));
	PE pe94_98(.x(x98),.w(w94_97),.acc(r94_97),.res(r94_98),.clk(clk),.wout(w94_98));
	PE pe94_99(.x(x99),.w(w94_98),.acc(r94_98),.res(r94_99),.clk(clk),.wout(w94_99));
	PE pe94_100(.x(x100),.w(w94_99),.acc(r94_99),.res(r94_100),.clk(clk),.wout(w94_100));
	PE pe94_101(.x(x101),.w(w94_100),.acc(r94_100),.res(r94_101),.clk(clk),.wout(w94_101));
	PE pe94_102(.x(x102),.w(w94_101),.acc(r94_101),.res(r94_102),.clk(clk),.wout(w94_102));
	PE pe94_103(.x(x103),.w(w94_102),.acc(r94_102),.res(r94_103),.clk(clk),.wout(w94_103));
	PE pe94_104(.x(x104),.w(w94_103),.acc(r94_103),.res(r94_104),.clk(clk),.wout(w94_104));
	PE pe94_105(.x(x105),.w(w94_104),.acc(r94_104),.res(r94_105),.clk(clk),.wout(w94_105));
	PE pe94_106(.x(x106),.w(w94_105),.acc(r94_105),.res(r94_106),.clk(clk),.wout(w94_106));
	PE pe94_107(.x(x107),.w(w94_106),.acc(r94_106),.res(r94_107),.clk(clk),.wout(w94_107));
	PE pe94_108(.x(x108),.w(w94_107),.acc(r94_107),.res(r94_108),.clk(clk),.wout(w94_108));
	PE pe94_109(.x(x109),.w(w94_108),.acc(r94_108),.res(r94_109),.clk(clk),.wout(w94_109));
	PE pe94_110(.x(x110),.w(w94_109),.acc(r94_109),.res(r94_110),.clk(clk),.wout(w94_110));
	PE pe94_111(.x(x111),.w(w94_110),.acc(r94_110),.res(r94_111),.clk(clk),.wout(w94_111));
	PE pe94_112(.x(x112),.w(w94_111),.acc(r94_111),.res(r94_112),.clk(clk),.wout(w94_112));
	PE pe94_113(.x(x113),.w(w94_112),.acc(r94_112),.res(r94_113),.clk(clk),.wout(w94_113));
	PE pe94_114(.x(x114),.w(w94_113),.acc(r94_113),.res(r94_114),.clk(clk),.wout(w94_114));
	PE pe94_115(.x(x115),.w(w94_114),.acc(r94_114),.res(r94_115),.clk(clk),.wout(w94_115));
	PE pe94_116(.x(x116),.w(w94_115),.acc(r94_115),.res(r94_116),.clk(clk),.wout(w94_116));
	PE pe94_117(.x(x117),.w(w94_116),.acc(r94_116),.res(r94_117),.clk(clk),.wout(w94_117));
	PE pe94_118(.x(x118),.w(w94_117),.acc(r94_117),.res(r94_118),.clk(clk),.wout(w94_118));
	PE pe94_119(.x(x119),.w(w94_118),.acc(r94_118),.res(r94_119),.clk(clk),.wout(w94_119));
	PE pe94_120(.x(x120),.w(w94_119),.acc(r94_119),.res(r94_120),.clk(clk),.wout(w94_120));
	PE pe94_121(.x(x121),.w(w94_120),.acc(r94_120),.res(r94_121),.clk(clk),.wout(w94_121));
	PE pe94_122(.x(x122),.w(w94_121),.acc(r94_121),.res(r94_122),.clk(clk),.wout(w94_122));
	PE pe94_123(.x(x123),.w(w94_122),.acc(r94_122),.res(r94_123),.clk(clk),.wout(w94_123));
	PE pe94_124(.x(x124),.w(w94_123),.acc(r94_123),.res(r94_124),.clk(clk),.wout(w94_124));
	PE pe94_125(.x(x125),.w(w94_124),.acc(r94_124),.res(r94_125),.clk(clk),.wout(w94_125));
	PE pe94_126(.x(x126),.w(w94_125),.acc(r94_125),.res(r94_126),.clk(clk),.wout(w94_126));
	PE pe94_127(.x(x127),.w(w94_126),.acc(r94_126),.res(result94),.clk(clk),.wout(weight94));

	PE pe95_0(.x(x0),.w(w95),.acc(32'h0),.res(r95_0),.clk(clk),.wout(w95_0));
	PE pe95_1(.x(x1),.w(w95_0),.acc(r95_0),.res(r95_1),.clk(clk),.wout(w95_1));
	PE pe95_2(.x(x2),.w(w95_1),.acc(r95_1),.res(r95_2),.clk(clk),.wout(w95_2));
	PE pe95_3(.x(x3),.w(w95_2),.acc(r95_2),.res(r95_3),.clk(clk),.wout(w95_3));
	PE pe95_4(.x(x4),.w(w95_3),.acc(r95_3),.res(r95_4),.clk(clk),.wout(w95_4));
	PE pe95_5(.x(x5),.w(w95_4),.acc(r95_4),.res(r95_5),.clk(clk),.wout(w95_5));
	PE pe95_6(.x(x6),.w(w95_5),.acc(r95_5),.res(r95_6),.clk(clk),.wout(w95_6));
	PE pe95_7(.x(x7),.w(w95_6),.acc(r95_6),.res(r95_7),.clk(clk),.wout(w95_7));
	PE pe95_8(.x(x8),.w(w95_7),.acc(r95_7),.res(r95_8),.clk(clk),.wout(w95_8));
	PE pe95_9(.x(x9),.w(w95_8),.acc(r95_8),.res(r95_9),.clk(clk),.wout(w95_9));
	PE pe95_10(.x(x10),.w(w95_9),.acc(r95_9),.res(r95_10),.clk(clk),.wout(w95_10));
	PE pe95_11(.x(x11),.w(w95_10),.acc(r95_10),.res(r95_11),.clk(clk),.wout(w95_11));
	PE pe95_12(.x(x12),.w(w95_11),.acc(r95_11),.res(r95_12),.clk(clk),.wout(w95_12));
	PE pe95_13(.x(x13),.w(w95_12),.acc(r95_12),.res(r95_13),.clk(clk),.wout(w95_13));
	PE pe95_14(.x(x14),.w(w95_13),.acc(r95_13),.res(r95_14),.clk(clk),.wout(w95_14));
	PE pe95_15(.x(x15),.w(w95_14),.acc(r95_14),.res(r95_15),.clk(clk),.wout(w95_15));
	PE pe95_16(.x(x16),.w(w95_15),.acc(r95_15),.res(r95_16),.clk(clk),.wout(w95_16));
	PE pe95_17(.x(x17),.w(w95_16),.acc(r95_16),.res(r95_17),.clk(clk),.wout(w95_17));
	PE pe95_18(.x(x18),.w(w95_17),.acc(r95_17),.res(r95_18),.clk(clk),.wout(w95_18));
	PE pe95_19(.x(x19),.w(w95_18),.acc(r95_18),.res(r95_19),.clk(clk),.wout(w95_19));
	PE pe95_20(.x(x20),.w(w95_19),.acc(r95_19),.res(r95_20),.clk(clk),.wout(w95_20));
	PE pe95_21(.x(x21),.w(w95_20),.acc(r95_20),.res(r95_21),.clk(clk),.wout(w95_21));
	PE pe95_22(.x(x22),.w(w95_21),.acc(r95_21),.res(r95_22),.clk(clk),.wout(w95_22));
	PE pe95_23(.x(x23),.w(w95_22),.acc(r95_22),.res(r95_23),.clk(clk),.wout(w95_23));
	PE pe95_24(.x(x24),.w(w95_23),.acc(r95_23),.res(r95_24),.clk(clk),.wout(w95_24));
	PE pe95_25(.x(x25),.w(w95_24),.acc(r95_24),.res(r95_25),.clk(clk),.wout(w95_25));
	PE pe95_26(.x(x26),.w(w95_25),.acc(r95_25),.res(r95_26),.clk(clk),.wout(w95_26));
	PE pe95_27(.x(x27),.w(w95_26),.acc(r95_26),.res(r95_27),.clk(clk),.wout(w95_27));
	PE pe95_28(.x(x28),.w(w95_27),.acc(r95_27),.res(r95_28),.clk(clk),.wout(w95_28));
	PE pe95_29(.x(x29),.w(w95_28),.acc(r95_28),.res(r95_29),.clk(clk),.wout(w95_29));
	PE pe95_30(.x(x30),.w(w95_29),.acc(r95_29),.res(r95_30),.clk(clk),.wout(w95_30));
	PE pe95_31(.x(x31),.w(w95_30),.acc(r95_30),.res(r95_31),.clk(clk),.wout(w95_31));
	PE pe95_32(.x(x32),.w(w95_31),.acc(r95_31),.res(r95_32),.clk(clk),.wout(w95_32));
	PE pe95_33(.x(x33),.w(w95_32),.acc(r95_32),.res(r95_33),.clk(clk),.wout(w95_33));
	PE pe95_34(.x(x34),.w(w95_33),.acc(r95_33),.res(r95_34),.clk(clk),.wout(w95_34));
	PE pe95_35(.x(x35),.w(w95_34),.acc(r95_34),.res(r95_35),.clk(clk),.wout(w95_35));
	PE pe95_36(.x(x36),.w(w95_35),.acc(r95_35),.res(r95_36),.clk(clk),.wout(w95_36));
	PE pe95_37(.x(x37),.w(w95_36),.acc(r95_36),.res(r95_37),.clk(clk),.wout(w95_37));
	PE pe95_38(.x(x38),.w(w95_37),.acc(r95_37),.res(r95_38),.clk(clk),.wout(w95_38));
	PE pe95_39(.x(x39),.w(w95_38),.acc(r95_38),.res(r95_39),.clk(clk),.wout(w95_39));
	PE pe95_40(.x(x40),.w(w95_39),.acc(r95_39),.res(r95_40),.clk(clk),.wout(w95_40));
	PE pe95_41(.x(x41),.w(w95_40),.acc(r95_40),.res(r95_41),.clk(clk),.wout(w95_41));
	PE pe95_42(.x(x42),.w(w95_41),.acc(r95_41),.res(r95_42),.clk(clk),.wout(w95_42));
	PE pe95_43(.x(x43),.w(w95_42),.acc(r95_42),.res(r95_43),.clk(clk),.wout(w95_43));
	PE pe95_44(.x(x44),.w(w95_43),.acc(r95_43),.res(r95_44),.clk(clk),.wout(w95_44));
	PE pe95_45(.x(x45),.w(w95_44),.acc(r95_44),.res(r95_45),.clk(clk),.wout(w95_45));
	PE pe95_46(.x(x46),.w(w95_45),.acc(r95_45),.res(r95_46),.clk(clk),.wout(w95_46));
	PE pe95_47(.x(x47),.w(w95_46),.acc(r95_46),.res(r95_47),.clk(clk),.wout(w95_47));
	PE pe95_48(.x(x48),.w(w95_47),.acc(r95_47),.res(r95_48),.clk(clk),.wout(w95_48));
	PE pe95_49(.x(x49),.w(w95_48),.acc(r95_48),.res(r95_49),.clk(clk),.wout(w95_49));
	PE pe95_50(.x(x50),.w(w95_49),.acc(r95_49),.res(r95_50),.clk(clk),.wout(w95_50));
	PE pe95_51(.x(x51),.w(w95_50),.acc(r95_50),.res(r95_51),.clk(clk),.wout(w95_51));
	PE pe95_52(.x(x52),.w(w95_51),.acc(r95_51),.res(r95_52),.clk(clk),.wout(w95_52));
	PE pe95_53(.x(x53),.w(w95_52),.acc(r95_52),.res(r95_53),.clk(clk),.wout(w95_53));
	PE pe95_54(.x(x54),.w(w95_53),.acc(r95_53),.res(r95_54),.clk(clk),.wout(w95_54));
	PE pe95_55(.x(x55),.w(w95_54),.acc(r95_54),.res(r95_55),.clk(clk),.wout(w95_55));
	PE pe95_56(.x(x56),.w(w95_55),.acc(r95_55),.res(r95_56),.clk(clk),.wout(w95_56));
	PE pe95_57(.x(x57),.w(w95_56),.acc(r95_56),.res(r95_57),.clk(clk),.wout(w95_57));
	PE pe95_58(.x(x58),.w(w95_57),.acc(r95_57),.res(r95_58),.clk(clk),.wout(w95_58));
	PE pe95_59(.x(x59),.w(w95_58),.acc(r95_58),.res(r95_59),.clk(clk),.wout(w95_59));
	PE pe95_60(.x(x60),.w(w95_59),.acc(r95_59),.res(r95_60),.clk(clk),.wout(w95_60));
	PE pe95_61(.x(x61),.w(w95_60),.acc(r95_60),.res(r95_61),.clk(clk),.wout(w95_61));
	PE pe95_62(.x(x62),.w(w95_61),.acc(r95_61),.res(r95_62),.clk(clk),.wout(w95_62));
	PE pe95_63(.x(x63),.w(w95_62),.acc(r95_62),.res(r95_63),.clk(clk),.wout(w95_63));
	PE pe95_64(.x(x64),.w(w95_63),.acc(r95_63),.res(r95_64),.clk(clk),.wout(w95_64));
	PE pe95_65(.x(x65),.w(w95_64),.acc(r95_64),.res(r95_65),.clk(clk),.wout(w95_65));
	PE pe95_66(.x(x66),.w(w95_65),.acc(r95_65),.res(r95_66),.clk(clk),.wout(w95_66));
	PE pe95_67(.x(x67),.w(w95_66),.acc(r95_66),.res(r95_67),.clk(clk),.wout(w95_67));
	PE pe95_68(.x(x68),.w(w95_67),.acc(r95_67),.res(r95_68),.clk(clk),.wout(w95_68));
	PE pe95_69(.x(x69),.w(w95_68),.acc(r95_68),.res(r95_69),.clk(clk),.wout(w95_69));
	PE pe95_70(.x(x70),.w(w95_69),.acc(r95_69),.res(r95_70),.clk(clk),.wout(w95_70));
	PE pe95_71(.x(x71),.w(w95_70),.acc(r95_70),.res(r95_71),.clk(clk),.wout(w95_71));
	PE pe95_72(.x(x72),.w(w95_71),.acc(r95_71),.res(r95_72),.clk(clk),.wout(w95_72));
	PE pe95_73(.x(x73),.w(w95_72),.acc(r95_72),.res(r95_73),.clk(clk),.wout(w95_73));
	PE pe95_74(.x(x74),.w(w95_73),.acc(r95_73),.res(r95_74),.clk(clk),.wout(w95_74));
	PE pe95_75(.x(x75),.w(w95_74),.acc(r95_74),.res(r95_75),.clk(clk),.wout(w95_75));
	PE pe95_76(.x(x76),.w(w95_75),.acc(r95_75),.res(r95_76),.clk(clk),.wout(w95_76));
	PE pe95_77(.x(x77),.w(w95_76),.acc(r95_76),.res(r95_77),.clk(clk),.wout(w95_77));
	PE pe95_78(.x(x78),.w(w95_77),.acc(r95_77),.res(r95_78),.clk(clk),.wout(w95_78));
	PE pe95_79(.x(x79),.w(w95_78),.acc(r95_78),.res(r95_79),.clk(clk),.wout(w95_79));
	PE pe95_80(.x(x80),.w(w95_79),.acc(r95_79),.res(r95_80),.clk(clk),.wout(w95_80));
	PE pe95_81(.x(x81),.w(w95_80),.acc(r95_80),.res(r95_81),.clk(clk),.wout(w95_81));
	PE pe95_82(.x(x82),.w(w95_81),.acc(r95_81),.res(r95_82),.clk(clk),.wout(w95_82));
	PE pe95_83(.x(x83),.w(w95_82),.acc(r95_82),.res(r95_83),.clk(clk),.wout(w95_83));
	PE pe95_84(.x(x84),.w(w95_83),.acc(r95_83),.res(r95_84),.clk(clk),.wout(w95_84));
	PE pe95_85(.x(x85),.w(w95_84),.acc(r95_84),.res(r95_85),.clk(clk),.wout(w95_85));
	PE pe95_86(.x(x86),.w(w95_85),.acc(r95_85),.res(r95_86),.clk(clk),.wout(w95_86));
	PE pe95_87(.x(x87),.w(w95_86),.acc(r95_86),.res(r95_87),.clk(clk),.wout(w95_87));
	PE pe95_88(.x(x88),.w(w95_87),.acc(r95_87),.res(r95_88),.clk(clk),.wout(w95_88));
	PE pe95_89(.x(x89),.w(w95_88),.acc(r95_88),.res(r95_89),.clk(clk),.wout(w95_89));
	PE pe95_90(.x(x90),.w(w95_89),.acc(r95_89),.res(r95_90),.clk(clk),.wout(w95_90));
	PE pe95_91(.x(x91),.w(w95_90),.acc(r95_90),.res(r95_91),.clk(clk),.wout(w95_91));
	PE pe95_92(.x(x92),.w(w95_91),.acc(r95_91),.res(r95_92),.clk(clk),.wout(w95_92));
	PE pe95_93(.x(x93),.w(w95_92),.acc(r95_92),.res(r95_93),.clk(clk),.wout(w95_93));
	PE pe95_94(.x(x94),.w(w95_93),.acc(r95_93),.res(r95_94),.clk(clk),.wout(w95_94));
	PE pe95_95(.x(x95),.w(w95_94),.acc(r95_94),.res(r95_95),.clk(clk),.wout(w95_95));
	PE pe95_96(.x(x96),.w(w95_95),.acc(r95_95),.res(r95_96),.clk(clk),.wout(w95_96));
	PE pe95_97(.x(x97),.w(w95_96),.acc(r95_96),.res(r95_97),.clk(clk),.wout(w95_97));
	PE pe95_98(.x(x98),.w(w95_97),.acc(r95_97),.res(r95_98),.clk(clk),.wout(w95_98));
	PE pe95_99(.x(x99),.w(w95_98),.acc(r95_98),.res(r95_99),.clk(clk),.wout(w95_99));
	PE pe95_100(.x(x100),.w(w95_99),.acc(r95_99),.res(r95_100),.clk(clk),.wout(w95_100));
	PE pe95_101(.x(x101),.w(w95_100),.acc(r95_100),.res(r95_101),.clk(clk),.wout(w95_101));
	PE pe95_102(.x(x102),.w(w95_101),.acc(r95_101),.res(r95_102),.clk(clk),.wout(w95_102));
	PE pe95_103(.x(x103),.w(w95_102),.acc(r95_102),.res(r95_103),.clk(clk),.wout(w95_103));
	PE pe95_104(.x(x104),.w(w95_103),.acc(r95_103),.res(r95_104),.clk(clk),.wout(w95_104));
	PE pe95_105(.x(x105),.w(w95_104),.acc(r95_104),.res(r95_105),.clk(clk),.wout(w95_105));
	PE pe95_106(.x(x106),.w(w95_105),.acc(r95_105),.res(r95_106),.clk(clk),.wout(w95_106));
	PE pe95_107(.x(x107),.w(w95_106),.acc(r95_106),.res(r95_107),.clk(clk),.wout(w95_107));
	PE pe95_108(.x(x108),.w(w95_107),.acc(r95_107),.res(r95_108),.clk(clk),.wout(w95_108));
	PE pe95_109(.x(x109),.w(w95_108),.acc(r95_108),.res(r95_109),.clk(clk),.wout(w95_109));
	PE pe95_110(.x(x110),.w(w95_109),.acc(r95_109),.res(r95_110),.clk(clk),.wout(w95_110));
	PE pe95_111(.x(x111),.w(w95_110),.acc(r95_110),.res(r95_111),.clk(clk),.wout(w95_111));
	PE pe95_112(.x(x112),.w(w95_111),.acc(r95_111),.res(r95_112),.clk(clk),.wout(w95_112));
	PE pe95_113(.x(x113),.w(w95_112),.acc(r95_112),.res(r95_113),.clk(clk),.wout(w95_113));
	PE pe95_114(.x(x114),.w(w95_113),.acc(r95_113),.res(r95_114),.clk(clk),.wout(w95_114));
	PE pe95_115(.x(x115),.w(w95_114),.acc(r95_114),.res(r95_115),.clk(clk),.wout(w95_115));
	PE pe95_116(.x(x116),.w(w95_115),.acc(r95_115),.res(r95_116),.clk(clk),.wout(w95_116));
	PE pe95_117(.x(x117),.w(w95_116),.acc(r95_116),.res(r95_117),.clk(clk),.wout(w95_117));
	PE pe95_118(.x(x118),.w(w95_117),.acc(r95_117),.res(r95_118),.clk(clk),.wout(w95_118));
	PE pe95_119(.x(x119),.w(w95_118),.acc(r95_118),.res(r95_119),.clk(clk),.wout(w95_119));
	PE pe95_120(.x(x120),.w(w95_119),.acc(r95_119),.res(r95_120),.clk(clk),.wout(w95_120));
	PE pe95_121(.x(x121),.w(w95_120),.acc(r95_120),.res(r95_121),.clk(clk),.wout(w95_121));
	PE pe95_122(.x(x122),.w(w95_121),.acc(r95_121),.res(r95_122),.clk(clk),.wout(w95_122));
	PE pe95_123(.x(x123),.w(w95_122),.acc(r95_122),.res(r95_123),.clk(clk),.wout(w95_123));
	PE pe95_124(.x(x124),.w(w95_123),.acc(r95_123),.res(r95_124),.clk(clk),.wout(w95_124));
	PE pe95_125(.x(x125),.w(w95_124),.acc(r95_124),.res(r95_125),.clk(clk),.wout(w95_125));
	PE pe95_126(.x(x126),.w(w95_125),.acc(r95_125),.res(r95_126),.clk(clk),.wout(w95_126));
	PE pe95_127(.x(x127),.w(w95_126),.acc(r95_126),.res(result95),.clk(clk),.wout(weight95));

	PE pe96_0(.x(x0),.w(w96),.acc(32'h0),.res(r96_0),.clk(clk),.wout(w96_0));
	PE pe96_1(.x(x1),.w(w96_0),.acc(r96_0),.res(r96_1),.clk(clk),.wout(w96_1));
	PE pe96_2(.x(x2),.w(w96_1),.acc(r96_1),.res(r96_2),.clk(clk),.wout(w96_2));
	PE pe96_3(.x(x3),.w(w96_2),.acc(r96_2),.res(r96_3),.clk(clk),.wout(w96_3));
	PE pe96_4(.x(x4),.w(w96_3),.acc(r96_3),.res(r96_4),.clk(clk),.wout(w96_4));
	PE pe96_5(.x(x5),.w(w96_4),.acc(r96_4),.res(r96_5),.clk(clk),.wout(w96_5));
	PE pe96_6(.x(x6),.w(w96_5),.acc(r96_5),.res(r96_6),.clk(clk),.wout(w96_6));
	PE pe96_7(.x(x7),.w(w96_6),.acc(r96_6),.res(r96_7),.clk(clk),.wout(w96_7));
	PE pe96_8(.x(x8),.w(w96_7),.acc(r96_7),.res(r96_8),.clk(clk),.wout(w96_8));
	PE pe96_9(.x(x9),.w(w96_8),.acc(r96_8),.res(r96_9),.clk(clk),.wout(w96_9));
	PE pe96_10(.x(x10),.w(w96_9),.acc(r96_9),.res(r96_10),.clk(clk),.wout(w96_10));
	PE pe96_11(.x(x11),.w(w96_10),.acc(r96_10),.res(r96_11),.clk(clk),.wout(w96_11));
	PE pe96_12(.x(x12),.w(w96_11),.acc(r96_11),.res(r96_12),.clk(clk),.wout(w96_12));
	PE pe96_13(.x(x13),.w(w96_12),.acc(r96_12),.res(r96_13),.clk(clk),.wout(w96_13));
	PE pe96_14(.x(x14),.w(w96_13),.acc(r96_13),.res(r96_14),.clk(clk),.wout(w96_14));
	PE pe96_15(.x(x15),.w(w96_14),.acc(r96_14),.res(r96_15),.clk(clk),.wout(w96_15));
	PE pe96_16(.x(x16),.w(w96_15),.acc(r96_15),.res(r96_16),.clk(clk),.wout(w96_16));
	PE pe96_17(.x(x17),.w(w96_16),.acc(r96_16),.res(r96_17),.clk(clk),.wout(w96_17));
	PE pe96_18(.x(x18),.w(w96_17),.acc(r96_17),.res(r96_18),.clk(clk),.wout(w96_18));
	PE pe96_19(.x(x19),.w(w96_18),.acc(r96_18),.res(r96_19),.clk(clk),.wout(w96_19));
	PE pe96_20(.x(x20),.w(w96_19),.acc(r96_19),.res(r96_20),.clk(clk),.wout(w96_20));
	PE pe96_21(.x(x21),.w(w96_20),.acc(r96_20),.res(r96_21),.clk(clk),.wout(w96_21));
	PE pe96_22(.x(x22),.w(w96_21),.acc(r96_21),.res(r96_22),.clk(clk),.wout(w96_22));
	PE pe96_23(.x(x23),.w(w96_22),.acc(r96_22),.res(r96_23),.clk(clk),.wout(w96_23));
	PE pe96_24(.x(x24),.w(w96_23),.acc(r96_23),.res(r96_24),.clk(clk),.wout(w96_24));
	PE pe96_25(.x(x25),.w(w96_24),.acc(r96_24),.res(r96_25),.clk(clk),.wout(w96_25));
	PE pe96_26(.x(x26),.w(w96_25),.acc(r96_25),.res(r96_26),.clk(clk),.wout(w96_26));
	PE pe96_27(.x(x27),.w(w96_26),.acc(r96_26),.res(r96_27),.clk(clk),.wout(w96_27));
	PE pe96_28(.x(x28),.w(w96_27),.acc(r96_27),.res(r96_28),.clk(clk),.wout(w96_28));
	PE pe96_29(.x(x29),.w(w96_28),.acc(r96_28),.res(r96_29),.clk(clk),.wout(w96_29));
	PE pe96_30(.x(x30),.w(w96_29),.acc(r96_29),.res(r96_30),.clk(clk),.wout(w96_30));
	PE pe96_31(.x(x31),.w(w96_30),.acc(r96_30),.res(r96_31),.clk(clk),.wout(w96_31));
	PE pe96_32(.x(x32),.w(w96_31),.acc(r96_31),.res(r96_32),.clk(clk),.wout(w96_32));
	PE pe96_33(.x(x33),.w(w96_32),.acc(r96_32),.res(r96_33),.clk(clk),.wout(w96_33));
	PE pe96_34(.x(x34),.w(w96_33),.acc(r96_33),.res(r96_34),.clk(clk),.wout(w96_34));
	PE pe96_35(.x(x35),.w(w96_34),.acc(r96_34),.res(r96_35),.clk(clk),.wout(w96_35));
	PE pe96_36(.x(x36),.w(w96_35),.acc(r96_35),.res(r96_36),.clk(clk),.wout(w96_36));
	PE pe96_37(.x(x37),.w(w96_36),.acc(r96_36),.res(r96_37),.clk(clk),.wout(w96_37));
	PE pe96_38(.x(x38),.w(w96_37),.acc(r96_37),.res(r96_38),.clk(clk),.wout(w96_38));
	PE pe96_39(.x(x39),.w(w96_38),.acc(r96_38),.res(r96_39),.clk(clk),.wout(w96_39));
	PE pe96_40(.x(x40),.w(w96_39),.acc(r96_39),.res(r96_40),.clk(clk),.wout(w96_40));
	PE pe96_41(.x(x41),.w(w96_40),.acc(r96_40),.res(r96_41),.clk(clk),.wout(w96_41));
	PE pe96_42(.x(x42),.w(w96_41),.acc(r96_41),.res(r96_42),.clk(clk),.wout(w96_42));
	PE pe96_43(.x(x43),.w(w96_42),.acc(r96_42),.res(r96_43),.clk(clk),.wout(w96_43));
	PE pe96_44(.x(x44),.w(w96_43),.acc(r96_43),.res(r96_44),.clk(clk),.wout(w96_44));
	PE pe96_45(.x(x45),.w(w96_44),.acc(r96_44),.res(r96_45),.clk(clk),.wout(w96_45));
	PE pe96_46(.x(x46),.w(w96_45),.acc(r96_45),.res(r96_46),.clk(clk),.wout(w96_46));
	PE pe96_47(.x(x47),.w(w96_46),.acc(r96_46),.res(r96_47),.clk(clk),.wout(w96_47));
	PE pe96_48(.x(x48),.w(w96_47),.acc(r96_47),.res(r96_48),.clk(clk),.wout(w96_48));
	PE pe96_49(.x(x49),.w(w96_48),.acc(r96_48),.res(r96_49),.clk(clk),.wout(w96_49));
	PE pe96_50(.x(x50),.w(w96_49),.acc(r96_49),.res(r96_50),.clk(clk),.wout(w96_50));
	PE pe96_51(.x(x51),.w(w96_50),.acc(r96_50),.res(r96_51),.clk(clk),.wout(w96_51));
	PE pe96_52(.x(x52),.w(w96_51),.acc(r96_51),.res(r96_52),.clk(clk),.wout(w96_52));
	PE pe96_53(.x(x53),.w(w96_52),.acc(r96_52),.res(r96_53),.clk(clk),.wout(w96_53));
	PE pe96_54(.x(x54),.w(w96_53),.acc(r96_53),.res(r96_54),.clk(clk),.wout(w96_54));
	PE pe96_55(.x(x55),.w(w96_54),.acc(r96_54),.res(r96_55),.clk(clk),.wout(w96_55));
	PE pe96_56(.x(x56),.w(w96_55),.acc(r96_55),.res(r96_56),.clk(clk),.wout(w96_56));
	PE pe96_57(.x(x57),.w(w96_56),.acc(r96_56),.res(r96_57),.clk(clk),.wout(w96_57));
	PE pe96_58(.x(x58),.w(w96_57),.acc(r96_57),.res(r96_58),.clk(clk),.wout(w96_58));
	PE pe96_59(.x(x59),.w(w96_58),.acc(r96_58),.res(r96_59),.clk(clk),.wout(w96_59));
	PE pe96_60(.x(x60),.w(w96_59),.acc(r96_59),.res(r96_60),.clk(clk),.wout(w96_60));
	PE pe96_61(.x(x61),.w(w96_60),.acc(r96_60),.res(r96_61),.clk(clk),.wout(w96_61));
	PE pe96_62(.x(x62),.w(w96_61),.acc(r96_61),.res(r96_62),.clk(clk),.wout(w96_62));
	PE pe96_63(.x(x63),.w(w96_62),.acc(r96_62),.res(r96_63),.clk(clk),.wout(w96_63));
	PE pe96_64(.x(x64),.w(w96_63),.acc(r96_63),.res(r96_64),.clk(clk),.wout(w96_64));
	PE pe96_65(.x(x65),.w(w96_64),.acc(r96_64),.res(r96_65),.clk(clk),.wout(w96_65));
	PE pe96_66(.x(x66),.w(w96_65),.acc(r96_65),.res(r96_66),.clk(clk),.wout(w96_66));
	PE pe96_67(.x(x67),.w(w96_66),.acc(r96_66),.res(r96_67),.clk(clk),.wout(w96_67));
	PE pe96_68(.x(x68),.w(w96_67),.acc(r96_67),.res(r96_68),.clk(clk),.wout(w96_68));
	PE pe96_69(.x(x69),.w(w96_68),.acc(r96_68),.res(r96_69),.clk(clk),.wout(w96_69));
	PE pe96_70(.x(x70),.w(w96_69),.acc(r96_69),.res(r96_70),.clk(clk),.wout(w96_70));
	PE pe96_71(.x(x71),.w(w96_70),.acc(r96_70),.res(r96_71),.clk(clk),.wout(w96_71));
	PE pe96_72(.x(x72),.w(w96_71),.acc(r96_71),.res(r96_72),.clk(clk),.wout(w96_72));
	PE pe96_73(.x(x73),.w(w96_72),.acc(r96_72),.res(r96_73),.clk(clk),.wout(w96_73));
	PE pe96_74(.x(x74),.w(w96_73),.acc(r96_73),.res(r96_74),.clk(clk),.wout(w96_74));
	PE pe96_75(.x(x75),.w(w96_74),.acc(r96_74),.res(r96_75),.clk(clk),.wout(w96_75));
	PE pe96_76(.x(x76),.w(w96_75),.acc(r96_75),.res(r96_76),.clk(clk),.wout(w96_76));
	PE pe96_77(.x(x77),.w(w96_76),.acc(r96_76),.res(r96_77),.clk(clk),.wout(w96_77));
	PE pe96_78(.x(x78),.w(w96_77),.acc(r96_77),.res(r96_78),.clk(clk),.wout(w96_78));
	PE pe96_79(.x(x79),.w(w96_78),.acc(r96_78),.res(r96_79),.clk(clk),.wout(w96_79));
	PE pe96_80(.x(x80),.w(w96_79),.acc(r96_79),.res(r96_80),.clk(clk),.wout(w96_80));
	PE pe96_81(.x(x81),.w(w96_80),.acc(r96_80),.res(r96_81),.clk(clk),.wout(w96_81));
	PE pe96_82(.x(x82),.w(w96_81),.acc(r96_81),.res(r96_82),.clk(clk),.wout(w96_82));
	PE pe96_83(.x(x83),.w(w96_82),.acc(r96_82),.res(r96_83),.clk(clk),.wout(w96_83));
	PE pe96_84(.x(x84),.w(w96_83),.acc(r96_83),.res(r96_84),.clk(clk),.wout(w96_84));
	PE pe96_85(.x(x85),.w(w96_84),.acc(r96_84),.res(r96_85),.clk(clk),.wout(w96_85));
	PE pe96_86(.x(x86),.w(w96_85),.acc(r96_85),.res(r96_86),.clk(clk),.wout(w96_86));
	PE pe96_87(.x(x87),.w(w96_86),.acc(r96_86),.res(r96_87),.clk(clk),.wout(w96_87));
	PE pe96_88(.x(x88),.w(w96_87),.acc(r96_87),.res(r96_88),.clk(clk),.wout(w96_88));
	PE pe96_89(.x(x89),.w(w96_88),.acc(r96_88),.res(r96_89),.clk(clk),.wout(w96_89));
	PE pe96_90(.x(x90),.w(w96_89),.acc(r96_89),.res(r96_90),.clk(clk),.wout(w96_90));
	PE pe96_91(.x(x91),.w(w96_90),.acc(r96_90),.res(r96_91),.clk(clk),.wout(w96_91));
	PE pe96_92(.x(x92),.w(w96_91),.acc(r96_91),.res(r96_92),.clk(clk),.wout(w96_92));
	PE pe96_93(.x(x93),.w(w96_92),.acc(r96_92),.res(r96_93),.clk(clk),.wout(w96_93));
	PE pe96_94(.x(x94),.w(w96_93),.acc(r96_93),.res(r96_94),.clk(clk),.wout(w96_94));
	PE pe96_95(.x(x95),.w(w96_94),.acc(r96_94),.res(r96_95),.clk(clk),.wout(w96_95));
	PE pe96_96(.x(x96),.w(w96_95),.acc(r96_95),.res(r96_96),.clk(clk),.wout(w96_96));
	PE pe96_97(.x(x97),.w(w96_96),.acc(r96_96),.res(r96_97),.clk(clk),.wout(w96_97));
	PE pe96_98(.x(x98),.w(w96_97),.acc(r96_97),.res(r96_98),.clk(clk),.wout(w96_98));
	PE pe96_99(.x(x99),.w(w96_98),.acc(r96_98),.res(r96_99),.clk(clk),.wout(w96_99));
	PE pe96_100(.x(x100),.w(w96_99),.acc(r96_99),.res(r96_100),.clk(clk),.wout(w96_100));
	PE pe96_101(.x(x101),.w(w96_100),.acc(r96_100),.res(r96_101),.clk(clk),.wout(w96_101));
	PE pe96_102(.x(x102),.w(w96_101),.acc(r96_101),.res(r96_102),.clk(clk),.wout(w96_102));
	PE pe96_103(.x(x103),.w(w96_102),.acc(r96_102),.res(r96_103),.clk(clk),.wout(w96_103));
	PE pe96_104(.x(x104),.w(w96_103),.acc(r96_103),.res(r96_104),.clk(clk),.wout(w96_104));
	PE pe96_105(.x(x105),.w(w96_104),.acc(r96_104),.res(r96_105),.clk(clk),.wout(w96_105));
	PE pe96_106(.x(x106),.w(w96_105),.acc(r96_105),.res(r96_106),.clk(clk),.wout(w96_106));
	PE pe96_107(.x(x107),.w(w96_106),.acc(r96_106),.res(r96_107),.clk(clk),.wout(w96_107));
	PE pe96_108(.x(x108),.w(w96_107),.acc(r96_107),.res(r96_108),.clk(clk),.wout(w96_108));
	PE pe96_109(.x(x109),.w(w96_108),.acc(r96_108),.res(r96_109),.clk(clk),.wout(w96_109));
	PE pe96_110(.x(x110),.w(w96_109),.acc(r96_109),.res(r96_110),.clk(clk),.wout(w96_110));
	PE pe96_111(.x(x111),.w(w96_110),.acc(r96_110),.res(r96_111),.clk(clk),.wout(w96_111));
	PE pe96_112(.x(x112),.w(w96_111),.acc(r96_111),.res(r96_112),.clk(clk),.wout(w96_112));
	PE pe96_113(.x(x113),.w(w96_112),.acc(r96_112),.res(r96_113),.clk(clk),.wout(w96_113));
	PE pe96_114(.x(x114),.w(w96_113),.acc(r96_113),.res(r96_114),.clk(clk),.wout(w96_114));
	PE pe96_115(.x(x115),.w(w96_114),.acc(r96_114),.res(r96_115),.clk(clk),.wout(w96_115));
	PE pe96_116(.x(x116),.w(w96_115),.acc(r96_115),.res(r96_116),.clk(clk),.wout(w96_116));
	PE pe96_117(.x(x117),.w(w96_116),.acc(r96_116),.res(r96_117),.clk(clk),.wout(w96_117));
	PE pe96_118(.x(x118),.w(w96_117),.acc(r96_117),.res(r96_118),.clk(clk),.wout(w96_118));
	PE pe96_119(.x(x119),.w(w96_118),.acc(r96_118),.res(r96_119),.clk(clk),.wout(w96_119));
	PE pe96_120(.x(x120),.w(w96_119),.acc(r96_119),.res(r96_120),.clk(clk),.wout(w96_120));
	PE pe96_121(.x(x121),.w(w96_120),.acc(r96_120),.res(r96_121),.clk(clk),.wout(w96_121));
	PE pe96_122(.x(x122),.w(w96_121),.acc(r96_121),.res(r96_122),.clk(clk),.wout(w96_122));
	PE pe96_123(.x(x123),.w(w96_122),.acc(r96_122),.res(r96_123),.clk(clk),.wout(w96_123));
	PE pe96_124(.x(x124),.w(w96_123),.acc(r96_123),.res(r96_124),.clk(clk),.wout(w96_124));
	PE pe96_125(.x(x125),.w(w96_124),.acc(r96_124),.res(r96_125),.clk(clk),.wout(w96_125));
	PE pe96_126(.x(x126),.w(w96_125),.acc(r96_125),.res(r96_126),.clk(clk),.wout(w96_126));
	PE pe96_127(.x(x127),.w(w96_126),.acc(r96_126),.res(result96),.clk(clk),.wout(weight96));

	PE pe97_0(.x(x0),.w(w97),.acc(32'h0),.res(r97_0),.clk(clk),.wout(w97_0));
	PE pe97_1(.x(x1),.w(w97_0),.acc(r97_0),.res(r97_1),.clk(clk),.wout(w97_1));
	PE pe97_2(.x(x2),.w(w97_1),.acc(r97_1),.res(r97_2),.clk(clk),.wout(w97_2));
	PE pe97_3(.x(x3),.w(w97_2),.acc(r97_2),.res(r97_3),.clk(clk),.wout(w97_3));
	PE pe97_4(.x(x4),.w(w97_3),.acc(r97_3),.res(r97_4),.clk(clk),.wout(w97_4));
	PE pe97_5(.x(x5),.w(w97_4),.acc(r97_4),.res(r97_5),.clk(clk),.wout(w97_5));
	PE pe97_6(.x(x6),.w(w97_5),.acc(r97_5),.res(r97_6),.clk(clk),.wout(w97_6));
	PE pe97_7(.x(x7),.w(w97_6),.acc(r97_6),.res(r97_7),.clk(clk),.wout(w97_7));
	PE pe97_8(.x(x8),.w(w97_7),.acc(r97_7),.res(r97_8),.clk(clk),.wout(w97_8));
	PE pe97_9(.x(x9),.w(w97_8),.acc(r97_8),.res(r97_9),.clk(clk),.wout(w97_9));
	PE pe97_10(.x(x10),.w(w97_9),.acc(r97_9),.res(r97_10),.clk(clk),.wout(w97_10));
	PE pe97_11(.x(x11),.w(w97_10),.acc(r97_10),.res(r97_11),.clk(clk),.wout(w97_11));
	PE pe97_12(.x(x12),.w(w97_11),.acc(r97_11),.res(r97_12),.clk(clk),.wout(w97_12));
	PE pe97_13(.x(x13),.w(w97_12),.acc(r97_12),.res(r97_13),.clk(clk),.wout(w97_13));
	PE pe97_14(.x(x14),.w(w97_13),.acc(r97_13),.res(r97_14),.clk(clk),.wout(w97_14));
	PE pe97_15(.x(x15),.w(w97_14),.acc(r97_14),.res(r97_15),.clk(clk),.wout(w97_15));
	PE pe97_16(.x(x16),.w(w97_15),.acc(r97_15),.res(r97_16),.clk(clk),.wout(w97_16));
	PE pe97_17(.x(x17),.w(w97_16),.acc(r97_16),.res(r97_17),.clk(clk),.wout(w97_17));
	PE pe97_18(.x(x18),.w(w97_17),.acc(r97_17),.res(r97_18),.clk(clk),.wout(w97_18));
	PE pe97_19(.x(x19),.w(w97_18),.acc(r97_18),.res(r97_19),.clk(clk),.wout(w97_19));
	PE pe97_20(.x(x20),.w(w97_19),.acc(r97_19),.res(r97_20),.clk(clk),.wout(w97_20));
	PE pe97_21(.x(x21),.w(w97_20),.acc(r97_20),.res(r97_21),.clk(clk),.wout(w97_21));
	PE pe97_22(.x(x22),.w(w97_21),.acc(r97_21),.res(r97_22),.clk(clk),.wout(w97_22));
	PE pe97_23(.x(x23),.w(w97_22),.acc(r97_22),.res(r97_23),.clk(clk),.wout(w97_23));
	PE pe97_24(.x(x24),.w(w97_23),.acc(r97_23),.res(r97_24),.clk(clk),.wout(w97_24));
	PE pe97_25(.x(x25),.w(w97_24),.acc(r97_24),.res(r97_25),.clk(clk),.wout(w97_25));
	PE pe97_26(.x(x26),.w(w97_25),.acc(r97_25),.res(r97_26),.clk(clk),.wout(w97_26));
	PE pe97_27(.x(x27),.w(w97_26),.acc(r97_26),.res(r97_27),.clk(clk),.wout(w97_27));
	PE pe97_28(.x(x28),.w(w97_27),.acc(r97_27),.res(r97_28),.clk(clk),.wout(w97_28));
	PE pe97_29(.x(x29),.w(w97_28),.acc(r97_28),.res(r97_29),.clk(clk),.wout(w97_29));
	PE pe97_30(.x(x30),.w(w97_29),.acc(r97_29),.res(r97_30),.clk(clk),.wout(w97_30));
	PE pe97_31(.x(x31),.w(w97_30),.acc(r97_30),.res(r97_31),.clk(clk),.wout(w97_31));
	PE pe97_32(.x(x32),.w(w97_31),.acc(r97_31),.res(r97_32),.clk(clk),.wout(w97_32));
	PE pe97_33(.x(x33),.w(w97_32),.acc(r97_32),.res(r97_33),.clk(clk),.wout(w97_33));
	PE pe97_34(.x(x34),.w(w97_33),.acc(r97_33),.res(r97_34),.clk(clk),.wout(w97_34));
	PE pe97_35(.x(x35),.w(w97_34),.acc(r97_34),.res(r97_35),.clk(clk),.wout(w97_35));
	PE pe97_36(.x(x36),.w(w97_35),.acc(r97_35),.res(r97_36),.clk(clk),.wout(w97_36));
	PE pe97_37(.x(x37),.w(w97_36),.acc(r97_36),.res(r97_37),.clk(clk),.wout(w97_37));
	PE pe97_38(.x(x38),.w(w97_37),.acc(r97_37),.res(r97_38),.clk(clk),.wout(w97_38));
	PE pe97_39(.x(x39),.w(w97_38),.acc(r97_38),.res(r97_39),.clk(clk),.wout(w97_39));
	PE pe97_40(.x(x40),.w(w97_39),.acc(r97_39),.res(r97_40),.clk(clk),.wout(w97_40));
	PE pe97_41(.x(x41),.w(w97_40),.acc(r97_40),.res(r97_41),.clk(clk),.wout(w97_41));
	PE pe97_42(.x(x42),.w(w97_41),.acc(r97_41),.res(r97_42),.clk(clk),.wout(w97_42));
	PE pe97_43(.x(x43),.w(w97_42),.acc(r97_42),.res(r97_43),.clk(clk),.wout(w97_43));
	PE pe97_44(.x(x44),.w(w97_43),.acc(r97_43),.res(r97_44),.clk(clk),.wout(w97_44));
	PE pe97_45(.x(x45),.w(w97_44),.acc(r97_44),.res(r97_45),.clk(clk),.wout(w97_45));
	PE pe97_46(.x(x46),.w(w97_45),.acc(r97_45),.res(r97_46),.clk(clk),.wout(w97_46));
	PE pe97_47(.x(x47),.w(w97_46),.acc(r97_46),.res(r97_47),.clk(clk),.wout(w97_47));
	PE pe97_48(.x(x48),.w(w97_47),.acc(r97_47),.res(r97_48),.clk(clk),.wout(w97_48));
	PE pe97_49(.x(x49),.w(w97_48),.acc(r97_48),.res(r97_49),.clk(clk),.wout(w97_49));
	PE pe97_50(.x(x50),.w(w97_49),.acc(r97_49),.res(r97_50),.clk(clk),.wout(w97_50));
	PE pe97_51(.x(x51),.w(w97_50),.acc(r97_50),.res(r97_51),.clk(clk),.wout(w97_51));
	PE pe97_52(.x(x52),.w(w97_51),.acc(r97_51),.res(r97_52),.clk(clk),.wout(w97_52));
	PE pe97_53(.x(x53),.w(w97_52),.acc(r97_52),.res(r97_53),.clk(clk),.wout(w97_53));
	PE pe97_54(.x(x54),.w(w97_53),.acc(r97_53),.res(r97_54),.clk(clk),.wout(w97_54));
	PE pe97_55(.x(x55),.w(w97_54),.acc(r97_54),.res(r97_55),.clk(clk),.wout(w97_55));
	PE pe97_56(.x(x56),.w(w97_55),.acc(r97_55),.res(r97_56),.clk(clk),.wout(w97_56));
	PE pe97_57(.x(x57),.w(w97_56),.acc(r97_56),.res(r97_57),.clk(clk),.wout(w97_57));
	PE pe97_58(.x(x58),.w(w97_57),.acc(r97_57),.res(r97_58),.clk(clk),.wout(w97_58));
	PE pe97_59(.x(x59),.w(w97_58),.acc(r97_58),.res(r97_59),.clk(clk),.wout(w97_59));
	PE pe97_60(.x(x60),.w(w97_59),.acc(r97_59),.res(r97_60),.clk(clk),.wout(w97_60));
	PE pe97_61(.x(x61),.w(w97_60),.acc(r97_60),.res(r97_61),.clk(clk),.wout(w97_61));
	PE pe97_62(.x(x62),.w(w97_61),.acc(r97_61),.res(r97_62),.clk(clk),.wout(w97_62));
	PE pe97_63(.x(x63),.w(w97_62),.acc(r97_62),.res(r97_63),.clk(clk),.wout(w97_63));
	PE pe97_64(.x(x64),.w(w97_63),.acc(r97_63),.res(r97_64),.clk(clk),.wout(w97_64));
	PE pe97_65(.x(x65),.w(w97_64),.acc(r97_64),.res(r97_65),.clk(clk),.wout(w97_65));
	PE pe97_66(.x(x66),.w(w97_65),.acc(r97_65),.res(r97_66),.clk(clk),.wout(w97_66));
	PE pe97_67(.x(x67),.w(w97_66),.acc(r97_66),.res(r97_67),.clk(clk),.wout(w97_67));
	PE pe97_68(.x(x68),.w(w97_67),.acc(r97_67),.res(r97_68),.clk(clk),.wout(w97_68));
	PE pe97_69(.x(x69),.w(w97_68),.acc(r97_68),.res(r97_69),.clk(clk),.wout(w97_69));
	PE pe97_70(.x(x70),.w(w97_69),.acc(r97_69),.res(r97_70),.clk(clk),.wout(w97_70));
	PE pe97_71(.x(x71),.w(w97_70),.acc(r97_70),.res(r97_71),.clk(clk),.wout(w97_71));
	PE pe97_72(.x(x72),.w(w97_71),.acc(r97_71),.res(r97_72),.clk(clk),.wout(w97_72));
	PE pe97_73(.x(x73),.w(w97_72),.acc(r97_72),.res(r97_73),.clk(clk),.wout(w97_73));
	PE pe97_74(.x(x74),.w(w97_73),.acc(r97_73),.res(r97_74),.clk(clk),.wout(w97_74));
	PE pe97_75(.x(x75),.w(w97_74),.acc(r97_74),.res(r97_75),.clk(clk),.wout(w97_75));
	PE pe97_76(.x(x76),.w(w97_75),.acc(r97_75),.res(r97_76),.clk(clk),.wout(w97_76));
	PE pe97_77(.x(x77),.w(w97_76),.acc(r97_76),.res(r97_77),.clk(clk),.wout(w97_77));
	PE pe97_78(.x(x78),.w(w97_77),.acc(r97_77),.res(r97_78),.clk(clk),.wout(w97_78));
	PE pe97_79(.x(x79),.w(w97_78),.acc(r97_78),.res(r97_79),.clk(clk),.wout(w97_79));
	PE pe97_80(.x(x80),.w(w97_79),.acc(r97_79),.res(r97_80),.clk(clk),.wout(w97_80));
	PE pe97_81(.x(x81),.w(w97_80),.acc(r97_80),.res(r97_81),.clk(clk),.wout(w97_81));
	PE pe97_82(.x(x82),.w(w97_81),.acc(r97_81),.res(r97_82),.clk(clk),.wout(w97_82));
	PE pe97_83(.x(x83),.w(w97_82),.acc(r97_82),.res(r97_83),.clk(clk),.wout(w97_83));
	PE pe97_84(.x(x84),.w(w97_83),.acc(r97_83),.res(r97_84),.clk(clk),.wout(w97_84));
	PE pe97_85(.x(x85),.w(w97_84),.acc(r97_84),.res(r97_85),.clk(clk),.wout(w97_85));
	PE pe97_86(.x(x86),.w(w97_85),.acc(r97_85),.res(r97_86),.clk(clk),.wout(w97_86));
	PE pe97_87(.x(x87),.w(w97_86),.acc(r97_86),.res(r97_87),.clk(clk),.wout(w97_87));
	PE pe97_88(.x(x88),.w(w97_87),.acc(r97_87),.res(r97_88),.clk(clk),.wout(w97_88));
	PE pe97_89(.x(x89),.w(w97_88),.acc(r97_88),.res(r97_89),.clk(clk),.wout(w97_89));
	PE pe97_90(.x(x90),.w(w97_89),.acc(r97_89),.res(r97_90),.clk(clk),.wout(w97_90));
	PE pe97_91(.x(x91),.w(w97_90),.acc(r97_90),.res(r97_91),.clk(clk),.wout(w97_91));
	PE pe97_92(.x(x92),.w(w97_91),.acc(r97_91),.res(r97_92),.clk(clk),.wout(w97_92));
	PE pe97_93(.x(x93),.w(w97_92),.acc(r97_92),.res(r97_93),.clk(clk),.wout(w97_93));
	PE pe97_94(.x(x94),.w(w97_93),.acc(r97_93),.res(r97_94),.clk(clk),.wout(w97_94));
	PE pe97_95(.x(x95),.w(w97_94),.acc(r97_94),.res(r97_95),.clk(clk),.wout(w97_95));
	PE pe97_96(.x(x96),.w(w97_95),.acc(r97_95),.res(r97_96),.clk(clk),.wout(w97_96));
	PE pe97_97(.x(x97),.w(w97_96),.acc(r97_96),.res(r97_97),.clk(clk),.wout(w97_97));
	PE pe97_98(.x(x98),.w(w97_97),.acc(r97_97),.res(r97_98),.clk(clk),.wout(w97_98));
	PE pe97_99(.x(x99),.w(w97_98),.acc(r97_98),.res(r97_99),.clk(clk),.wout(w97_99));
	PE pe97_100(.x(x100),.w(w97_99),.acc(r97_99),.res(r97_100),.clk(clk),.wout(w97_100));
	PE pe97_101(.x(x101),.w(w97_100),.acc(r97_100),.res(r97_101),.clk(clk),.wout(w97_101));
	PE pe97_102(.x(x102),.w(w97_101),.acc(r97_101),.res(r97_102),.clk(clk),.wout(w97_102));
	PE pe97_103(.x(x103),.w(w97_102),.acc(r97_102),.res(r97_103),.clk(clk),.wout(w97_103));
	PE pe97_104(.x(x104),.w(w97_103),.acc(r97_103),.res(r97_104),.clk(clk),.wout(w97_104));
	PE pe97_105(.x(x105),.w(w97_104),.acc(r97_104),.res(r97_105),.clk(clk),.wout(w97_105));
	PE pe97_106(.x(x106),.w(w97_105),.acc(r97_105),.res(r97_106),.clk(clk),.wout(w97_106));
	PE pe97_107(.x(x107),.w(w97_106),.acc(r97_106),.res(r97_107),.clk(clk),.wout(w97_107));
	PE pe97_108(.x(x108),.w(w97_107),.acc(r97_107),.res(r97_108),.clk(clk),.wout(w97_108));
	PE pe97_109(.x(x109),.w(w97_108),.acc(r97_108),.res(r97_109),.clk(clk),.wout(w97_109));
	PE pe97_110(.x(x110),.w(w97_109),.acc(r97_109),.res(r97_110),.clk(clk),.wout(w97_110));
	PE pe97_111(.x(x111),.w(w97_110),.acc(r97_110),.res(r97_111),.clk(clk),.wout(w97_111));
	PE pe97_112(.x(x112),.w(w97_111),.acc(r97_111),.res(r97_112),.clk(clk),.wout(w97_112));
	PE pe97_113(.x(x113),.w(w97_112),.acc(r97_112),.res(r97_113),.clk(clk),.wout(w97_113));
	PE pe97_114(.x(x114),.w(w97_113),.acc(r97_113),.res(r97_114),.clk(clk),.wout(w97_114));
	PE pe97_115(.x(x115),.w(w97_114),.acc(r97_114),.res(r97_115),.clk(clk),.wout(w97_115));
	PE pe97_116(.x(x116),.w(w97_115),.acc(r97_115),.res(r97_116),.clk(clk),.wout(w97_116));
	PE pe97_117(.x(x117),.w(w97_116),.acc(r97_116),.res(r97_117),.clk(clk),.wout(w97_117));
	PE pe97_118(.x(x118),.w(w97_117),.acc(r97_117),.res(r97_118),.clk(clk),.wout(w97_118));
	PE pe97_119(.x(x119),.w(w97_118),.acc(r97_118),.res(r97_119),.clk(clk),.wout(w97_119));
	PE pe97_120(.x(x120),.w(w97_119),.acc(r97_119),.res(r97_120),.clk(clk),.wout(w97_120));
	PE pe97_121(.x(x121),.w(w97_120),.acc(r97_120),.res(r97_121),.clk(clk),.wout(w97_121));
	PE pe97_122(.x(x122),.w(w97_121),.acc(r97_121),.res(r97_122),.clk(clk),.wout(w97_122));
	PE pe97_123(.x(x123),.w(w97_122),.acc(r97_122),.res(r97_123),.clk(clk),.wout(w97_123));
	PE pe97_124(.x(x124),.w(w97_123),.acc(r97_123),.res(r97_124),.clk(clk),.wout(w97_124));
	PE pe97_125(.x(x125),.w(w97_124),.acc(r97_124),.res(r97_125),.clk(clk),.wout(w97_125));
	PE pe97_126(.x(x126),.w(w97_125),.acc(r97_125),.res(r97_126),.clk(clk),.wout(w97_126));
	PE pe97_127(.x(x127),.w(w97_126),.acc(r97_126),.res(result97),.clk(clk),.wout(weight97));

	PE pe98_0(.x(x0),.w(w98),.acc(32'h0),.res(r98_0),.clk(clk),.wout(w98_0));
	PE pe98_1(.x(x1),.w(w98_0),.acc(r98_0),.res(r98_1),.clk(clk),.wout(w98_1));
	PE pe98_2(.x(x2),.w(w98_1),.acc(r98_1),.res(r98_2),.clk(clk),.wout(w98_2));
	PE pe98_3(.x(x3),.w(w98_2),.acc(r98_2),.res(r98_3),.clk(clk),.wout(w98_3));
	PE pe98_4(.x(x4),.w(w98_3),.acc(r98_3),.res(r98_4),.clk(clk),.wout(w98_4));
	PE pe98_5(.x(x5),.w(w98_4),.acc(r98_4),.res(r98_5),.clk(clk),.wout(w98_5));
	PE pe98_6(.x(x6),.w(w98_5),.acc(r98_5),.res(r98_6),.clk(clk),.wout(w98_6));
	PE pe98_7(.x(x7),.w(w98_6),.acc(r98_6),.res(r98_7),.clk(clk),.wout(w98_7));
	PE pe98_8(.x(x8),.w(w98_7),.acc(r98_7),.res(r98_8),.clk(clk),.wout(w98_8));
	PE pe98_9(.x(x9),.w(w98_8),.acc(r98_8),.res(r98_9),.clk(clk),.wout(w98_9));
	PE pe98_10(.x(x10),.w(w98_9),.acc(r98_9),.res(r98_10),.clk(clk),.wout(w98_10));
	PE pe98_11(.x(x11),.w(w98_10),.acc(r98_10),.res(r98_11),.clk(clk),.wout(w98_11));
	PE pe98_12(.x(x12),.w(w98_11),.acc(r98_11),.res(r98_12),.clk(clk),.wout(w98_12));
	PE pe98_13(.x(x13),.w(w98_12),.acc(r98_12),.res(r98_13),.clk(clk),.wout(w98_13));
	PE pe98_14(.x(x14),.w(w98_13),.acc(r98_13),.res(r98_14),.clk(clk),.wout(w98_14));
	PE pe98_15(.x(x15),.w(w98_14),.acc(r98_14),.res(r98_15),.clk(clk),.wout(w98_15));
	PE pe98_16(.x(x16),.w(w98_15),.acc(r98_15),.res(r98_16),.clk(clk),.wout(w98_16));
	PE pe98_17(.x(x17),.w(w98_16),.acc(r98_16),.res(r98_17),.clk(clk),.wout(w98_17));
	PE pe98_18(.x(x18),.w(w98_17),.acc(r98_17),.res(r98_18),.clk(clk),.wout(w98_18));
	PE pe98_19(.x(x19),.w(w98_18),.acc(r98_18),.res(r98_19),.clk(clk),.wout(w98_19));
	PE pe98_20(.x(x20),.w(w98_19),.acc(r98_19),.res(r98_20),.clk(clk),.wout(w98_20));
	PE pe98_21(.x(x21),.w(w98_20),.acc(r98_20),.res(r98_21),.clk(clk),.wout(w98_21));
	PE pe98_22(.x(x22),.w(w98_21),.acc(r98_21),.res(r98_22),.clk(clk),.wout(w98_22));
	PE pe98_23(.x(x23),.w(w98_22),.acc(r98_22),.res(r98_23),.clk(clk),.wout(w98_23));
	PE pe98_24(.x(x24),.w(w98_23),.acc(r98_23),.res(r98_24),.clk(clk),.wout(w98_24));
	PE pe98_25(.x(x25),.w(w98_24),.acc(r98_24),.res(r98_25),.clk(clk),.wout(w98_25));
	PE pe98_26(.x(x26),.w(w98_25),.acc(r98_25),.res(r98_26),.clk(clk),.wout(w98_26));
	PE pe98_27(.x(x27),.w(w98_26),.acc(r98_26),.res(r98_27),.clk(clk),.wout(w98_27));
	PE pe98_28(.x(x28),.w(w98_27),.acc(r98_27),.res(r98_28),.clk(clk),.wout(w98_28));
	PE pe98_29(.x(x29),.w(w98_28),.acc(r98_28),.res(r98_29),.clk(clk),.wout(w98_29));
	PE pe98_30(.x(x30),.w(w98_29),.acc(r98_29),.res(r98_30),.clk(clk),.wout(w98_30));
	PE pe98_31(.x(x31),.w(w98_30),.acc(r98_30),.res(r98_31),.clk(clk),.wout(w98_31));
	PE pe98_32(.x(x32),.w(w98_31),.acc(r98_31),.res(r98_32),.clk(clk),.wout(w98_32));
	PE pe98_33(.x(x33),.w(w98_32),.acc(r98_32),.res(r98_33),.clk(clk),.wout(w98_33));
	PE pe98_34(.x(x34),.w(w98_33),.acc(r98_33),.res(r98_34),.clk(clk),.wout(w98_34));
	PE pe98_35(.x(x35),.w(w98_34),.acc(r98_34),.res(r98_35),.clk(clk),.wout(w98_35));
	PE pe98_36(.x(x36),.w(w98_35),.acc(r98_35),.res(r98_36),.clk(clk),.wout(w98_36));
	PE pe98_37(.x(x37),.w(w98_36),.acc(r98_36),.res(r98_37),.clk(clk),.wout(w98_37));
	PE pe98_38(.x(x38),.w(w98_37),.acc(r98_37),.res(r98_38),.clk(clk),.wout(w98_38));
	PE pe98_39(.x(x39),.w(w98_38),.acc(r98_38),.res(r98_39),.clk(clk),.wout(w98_39));
	PE pe98_40(.x(x40),.w(w98_39),.acc(r98_39),.res(r98_40),.clk(clk),.wout(w98_40));
	PE pe98_41(.x(x41),.w(w98_40),.acc(r98_40),.res(r98_41),.clk(clk),.wout(w98_41));
	PE pe98_42(.x(x42),.w(w98_41),.acc(r98_41),.res(r98_42),.clk(clk),.wout(w98_42));
	PE pe98_43(.x(x43),.w(w98_42),.acc(r98_42),.res(r98_43),.clk(clk),.wout(w98_43));
	PE pe98_44(.x(x44),.w(w98_43),.acc(r98_43),.res(r98_44),.clk(clk),.wout(w98_44));
	PE pe98_45(.x(x45),.w(w98_44),.acc(r98_44),.res(r98_45),.clk(clk),.wout(w98_45));
	PE pe98_46(.x(x46),.w(w98_45),.acc(r98_45),.res(r98_46),.clk(clk),.wout(w98_46));
	PE pe98_47(.x(x47),.w(w98_46),.acc(r98_46),.res(r98_47),.clk(clk),.wout(w98_47));
	PE pe98_48(.x(x48),.w(w98_47),.acc(r98_47),.res(r98_48),.clk(clk),.wout(w98_48));
	PE pe98_49(.x(x49),.w(w98_48),.acc(r98_48),.res(r98_49),.clk(clk),.wout(w98_49));
	PE pe98_50(.x(x50),.w(w98_49),.acc(r98_49),.res(r98_50),.clk(clk),.wout(w98_50));
	PE pe98_51(.x(x51),.w(w98_50),.acc(r98_50),.res(r98_51),.clk(clk),.wout(w98_51));
	PE pe98_52(.x(x52),.w(w98_51),.acc(r98_51),.res(r98_52),.clk(clk),.wout(w98_52));
	PE pe98_53(.x(x53),.w(w98_52),.acc(r98_52),.res(r98_53),.clk(clk),.wout(w98_53));
	PE pe98_54(.x(x54),.w(w98_53),.acc(r98_53),.res(r98_54),.clk(clk),.wout(w98_54));
	PE pe98_55(.x(x55),.w(w98_54),.acc(r98_54),.res(r98_55),.clk(clk),.wout(w98_55));
	PE pe98_56(.x(x56),.w(w98_55),.acc(r98_55),.res(r98_56),.clk(clk),.wout(w98_56));
	PE pe98_57(.x(x57),.w(w98_56),.acc(r98_56),.res(r98_57),.clk(clk),.wout(w98_57));
	PE pe98_58(.x(x58),.w(w98_57),.acc(r98_57),.res(r98_58),.clk(clk),.wout(w98_58));
	PE pe98_59(.x(x59),.w(w98_58),.acc(r98_58),.res(r98_59),.clk(clk),.wout(w98_59));
	PE pe98_60(.x(x60),.w(w98_59),.acc(r98_59),.res(r98_60),.clk(clk),.wout(w98_60));
	PE pe98_61(.x(x61),.w(w98_60),.acc(r98_60),.res(r98_61),.clk(clk),.wout(w98_61));
	PE pe98_62(.x(x62),.w(w98_61),.acc(r98_61),.res(r98_62),.clk(clk),.wout(w98_62));
	PE pe98_63(.x(x63),.w(w98_62),.acc(r98_62),.res(r98_63),.clk(clk),.wout(w98_63));
	PE pe98_64(.x(x64),.w(w98_63),.acc(r98_63),.res(r98_64),.clk(clk),.wout(w98_64));
	PE pe98_65(.x(x65),.w(w98_64),.acc(r98_64),.res(r98_65),.clk(clk),.wout(w98_65));
	PE pe98_66(.x(x66),.w(w98_65),.acc(r98_65),.res(r98_66),.clk(clk),.wout(w98_66));
	PE pe98_67(.x(x67),.w(w98_66),.acc(r98_66),.res(r98_67),.clk(clk),.wout(w98_67));
	PE pe98_68(.x(x68),.w(w98_67),.acc(r98_67),.res(r98_68),.clk(clk),.wout(w98_68));
	PE pe98_69(.x(x69),.w(w98_68),.acc(r98_68),.res(r98_69),.clk(clk),.wout(w98_69));
	PE pe98_70(.x(x70),.w(w98_69),.acc(r98_69),.res(r98_70),.clk(clk),.wout(w98_70));
	PE pe98_71(.x(x71),.w(w98_70),.acc(r98_70),.res(r98_71),.clk(clk),.wout(w98_71));
	PE pe98_72(.x(x72),.w(w98_71),.acc(r98_71),.res(r98_72),.clk(clk),.wout(w98_72));
	PE pe98_73(.x(x73),.w(w98_72),.acc(r98_72),.res(r98_73),.clk(clk),.wout(w98_73));
	PE pe98_74(.x(x74),.w(w98_73),.acc(r98_73),.res(r98_74),.clk(clk),.wout(w98_74));
	PE pe98_75(.x(x75),.w(w98_74),.acc(r98_74),.res(r98_75),.clk(clk),.wout(w98_75));
	PE pe98_76(.x(x76),.w(w98_75),.acc(r98_75),.res(r98_76),.clk(clk),.wout(w98_76));
	PE pe98_77(.x(x77),.w(w98_76),.acc(r98_76),.res(r98_77),.clk(clk),.wout(w98_77));
	PE pe98_78(.x(x78),.w(w98_77),.acc(r98_77),.res(r98_78),.clk(clk),.wout(w98_78));
	PE pe98_79(.x(x79),.w(w98_78),.acc(r98_78),.res(r98_79),.clk(clk),.wout(w98_79));
	PE pe98_80(.x(x80),.w(w98_79),.acc(r98_79),.res(r98_80),.clk(clk),.wout(w98_80));
	PE pe98_81(.x(x81),.w(w98_80),.acc(r98_80),.res(r98_81),.clk(clk),.wout(w98_81));
	PE pe98_82(.x(x82),.w(w98_81),.acc(r98_81),.res(r98_82),.clk(clk),.wout(w98_82));
	PE pe98_83(.x(x83),.w(w98_82),.acc(r98_82),.res(r98_83),.clk(clk),.wout(w98_83));
	PE pe98_84(.x(x84),.w(w98_83),.acc(r98_83),.res(r98_84),.clk(clk),.wout(w98_84));
	PE pe98_85(.x(x85),.w(w98_84),.acc(r98_84),.res(r98_85),.clk(clk),.wout(w98_85));
	PE pe98_86(.x(x86),.w(w98_85),.acc(r98_85),.res(r98_86),.clk(clk),.wout(w98_86));
	PE pe98_87(.x(x87),.w(w98_86),.acc(r98_86),.res(r98_87),.clk(clk),.wout(w98_87));
	PE pe98_88(.x(x88),.w(w98_87),.acc(r98_87),.res(r98_88),.clk(clk),.wout(w98_88));
	PE pe98_89(.x(x89),.w(w98_88),.acc(r98_88),.res(r98_89),.clk(clk),.wout(w98_89));
	PE pe98_90(.x(x90),.w(w98_89),.acc(r98_89),.res(r98_90),.clk(clk),.wout(w98_90));
	PE pe98_91(.x(x91),.w(w98_90),.acc(r98_90),.res(r98_91),.clk(clk),.wout(w98_91));
	PE pe98_92(.x(x92),.w(w98_91),.acc(r98_91),.res(r98_92),.clk(clk),.wout(w98_92));
	PE pe98_93(.x(x93),.w(w98_92),.acc(r98_92),.res(r98_93),.clk(clk),.wout(w98_93));
	PE pe98_94(.x(x94),.w(w98_93),.acc(r98_93),.res(r98_94),.clk(clk),.wout(w98_94));
	PE pe98_95(.x(x95),.w(w98_94),.acc(r98_94),.res(r98_95),.clk(clk),.wout(w98_95));
	PE pe98_96(.x(x96),.w(w98_95),.acc(r98_95),.res(r98_96),.clk(clk),.wout(w98_96));
	PE pe98_97(.x(x97),.w(w98_96),.acc(r98_96),.res(r98_97),.clk(clk),.wout(w98_97));
	PE pe98_98(.x(x98),.w(w98_97),.acc(r98_97),.res(r98_98),.clk(clk),.wout(w98_98));
	PE pe98_99(.x(x99),.w(w98_98),.acc(r98_98),.res(r98_99),.clk(clk),.wout(w98_99));
	PE pe98_100(.x(x100),.w(w98_99),.acc(r98_99),.res(r98_100),.clk(clk),.wout(w98_100));
	PE pe98_101(.x(x101),.w(w98_100),.acc(r98_100),.res(r98_101),.clk(clk),.wout(w98_101));
	PE pe98_102(.x(x102),.w(w98_101),.acc(r98_101),.res(r98_102),.clk(clk),.wout(w98_102));
	PE pe98_103(.x(x103),.w(w98_102),.acc(r98_102),.res(r98_103),.clk(clk),.wout(w98_103));
	PE pe98_104(.x(x104),.w(w98_103),.acc(r98_103),.res(r98_104),.clk(clk),.wout(w98_104));
	PE pe98_105(.x(x105),.w(w98_104),.acc(r98_104),.res(r98_105),.clk(clk),.wout(w98_105));
	PE pe98_106(.x(x106),.w(w98_105),.acc(r98_105),.res(r98_106),.clk(clk),.wout(w98_106));
	PE pe98_107(.x(x107),.w(w98_106),.acc(r98_106),.res(r98_107),.clk(clk),.wout(w98_107));
	PE pe98_108(.x(x108),.w(w98_107),.acc(r98_107),.res(r98_108),.clk(clk),.wout(w98_108));
	PE pe98_109(.x(x109),.w(w98_108),.acc(r98_108),.res(r98_109),.clk(clk),.wout(w98_109));
	PE pe98_110(.x(x110),.w(w98_109),.acc(r98_109),.res(r98_110),.clk(clk),.wout(w98_110));
	PE pe98_111(.x(x111),.w(w98_110),.acc(r98_110),.res(r98_111),.clk(clk),.wout(w98_111));
	PE pe98_112(.x(x112),.w(w98_111),.acc(r98_111),.res(r98_112),.clk(clk),.wout(w98_112));
	PE pe98_113(.x(x113),.w(w98_112),.acc(r98_112),.res(r98_113),.clk(clk),.wout(w98_113));
	PE pe98_114(.x(x114),.w(w98_113),.acc(r98_113),.res(r98_114),.clk(clk),.wout(w98_114));
	PE pe98_115(.x(x115),.w(w98_114),.acc(r98_114),.res(r98_115),.clk(clk),.wout(w98_115));
	PE pe98_116(.x(x116),.w(w98_115),.acc(r98_115),.res(r98_116),.clk(clk),.wout(w98_116));
	PE pe98_117(.x(x117),.w(w98_116),.acc(r98_116),.res(r98_117),.clk(clk),.wout(w98_117));
	PE pe98_118(.x(x118),.w(w98_117),.acc(r98_117),.res(r98_118),.clk(clk),.wout(w98_118));
	PE pe98_119(.x(x119),.w(w98_118),.acc(r98_118),.res(r98_119),.clk(clk),.wout(w98_119));
	PE pe98_120(.x(x120),.w(w98_119),.acc(r98_119),.res(r98_120),.clk(clk),.wout(w98_120));
	PE pe98_121(.x(x121),.w(w98_120),.acc(r98_120),.res(r98_121),.clk(clk),.wout(w98_121));
	PE pe98_122(.x(x122),.w(w98_121),.acc(r98_121),.res(r98_122),.clk(clk),.wout(w98_122));
	PE pe98_123(.x(x123),.w(w98_122),.acc(r98_122),.res(r98_123),.clk(clk),.wout(w98_123));
	PE pe98_124(.x(x124),.w(w98_123),.acc(r98_123),.res(r98_124),.clk(clk),.wout(w98_124));
	PE pe98_125(.x(x125),.w(w98_124),.acc(r98_124),.res(r98_125),.clk(clk),.wout(w98_125));
	PE pe98_126(.x(x126),.w(w98_125),.acc(r98_125),.res(r98_126),.clk(clk),.wout(w98_126));
	PE pe98_127(.x(x127),.w(w98_126),.acc(r98_126),.res(result98),.clk(clk),.wout(weight98));

	PE pe99_0(.x(x0),.w(w99),.acc(32'h0),.res(r99_0),.clk(clk),.wout(w99_0));
	PE pe99_1(.x(x1),.w(w99_0),.acc(r99_0),.res(r99_1),.clk(clk),.wout(w99_1));
	PE pe99_2(.x(x2),.w(w99_1),.acc(r99_1),.res(r99_2),.clk(clk),.wout(w99_2));
	PE pe99_3(.x(x3),.w(w99_2),.acc(r99_2),.res(r99_3),.clk(clk),.wout(w99_3));
	PE pe99_4(.x(x4),.w(w99_3),.acc(r99_3),.res(r99_4),.clk(clk),.wout(w99_4));
	PE pe99_5(.x(x5),.w(w99_4),.acc(r99_4),.res(r99_5),.clk(clk),.wout(w99_5));
	PE pe99_6(.x(x6),.w(w99_5),.acc(r99_5),.res(r99_6),.clk(clk),.wout(w99_6));
	PE pe99_7(.x(x7),.w(w99_6),.acc(r99_6),.res(r99_7),.clk(clk),.wout(w99_7));
	PE pe99_8(.x(x8),.w(w99_7),.acc(r99_7),.res(r99_8),.clk(clk),.wout(w99_8));
	PE pe99_9(.x(x9),.w(w99_8),.acc(r99_8),.res(r99_9),.clk(clk),.wout(w99_9));
	PE pe99_10(.x(x10),.w(w99_9),.acc(r99_9),.res(r99_10),.clk(clk),.wout(w99_10));
	PE pe99_11(.x(x11),.w(w99_10),.acc(r99_10),.res(r99_11),.clk(clk),.wout(w99_11));
	PE pe99_12(.x(x12),.w(w99_11),.acc(r99_11),.res(r99_12),.clk(clk),.wout(w99_12));
	PE pe99_13(.x(x13),.w(w99_12),.acc(r99_12),.res(r99_13),.clk(clk),.wout(w99_13));
	PE pe99_14(.x(x14),.w(w99_13),.acc(r99_13),.res(r99_14),.clk(clk),.wout(w99_14));
	PE pe99_15(.x(x15),.w(w99_14),.acc(r99_14),.res(r99_15),.clk(clk),.wout(w99_15));
	PE pe99_16(.x(x16),.w(w99_15),.acc(r99_15),.res(r99_16),.clk(clk),.wout(w99_16));
	PE pe99_17(.x(x17),.w(w99_16),.acc(r99_16),.res(r99_17),.clk(clk),.wout(w99_17));
	PE pe99_18(.x(x18),.w(w99_17),.acc(r99_17),.res(r99_18),.clk(clk),.wout(w99_18));
	PE pe99_19(.x(x19),.w(w99_18),.acc(r99_18),.res(r99_19),.clk(clk),.wout(w99_19));
	PE pe99_20(.x(x20),.w(w99_19),.acc(r99_19),.res(r99_20),.clk(clk),.wout(w99_20));
	PE pe99_21(.x(x21),.w(w99_20),.acc(r99_20),.res(r99_21),.clk(clk),.wout(w99_21));
	PE pe99_22(.x(x22),.w(w99_21),.acc(r99_21),.res(r99_22),.clk(clk),.wout(w99_22));
	PE pe99_23(.x(x23),.w(w99_22),.acc(r99_22),.res(r99_23),.clk(clk),.wout(w99_23));
	PE pe99_24(.x(x24),.w(w99_23),.acc(r99_23),.res(r99_24),.clk(clk),.wout(w99_24));
	PE pe99_25(.x(x25),.w(w99_24),.acc(r99_24),.res(r99_25),.clk(clk),.wout(w99_25));
	PE pe99_26(.x(x26),.w(w99_25),.acc(r99_25),.res(r99_26),.clk(clk),.wout(w99_26));
	PE pe99_27(.x(x27),.w(w99_26),.acc(r99_26),.res(r99_27),.clk(clk),.wout(w99_27));
	PE pe99_28(.x(x28),.w(w99_27),.acc(r99_27),.res(r99_28),.clk(clk),.wout(w99_28));
	PE pe99_29(.x(x29),.w(w99_28),.acc(r99_28),.res(r99_29),.clk(clk),.wout(w99_29));
	PE pe99_30(.x(x30),.w(w99_29),.acc(r99_29),.res(r99_30),.clk(clk),.wout(w99_30));
	PE pe99_31(.x(x31),.w(w99_30),.acc(r99_30),.res(r99_31),.clk(clk),.wout(w99_31));
	PE pe99_32(.x(x32),.w(w99_31),.acc(r99_31),.res(r99_32),.clk(clk),.wout(w99_32));
	PE pe99_33(.x(x33),.w(w99_32),.acc(r99_32),.res(r99_33),.clk(clk),.wout(w99_33));
	PE pe99_34(.x(x34),.w(w99_33),.acc(r99_33),.res(r99_34),.clk(clk),.wout(w99_34));
	PE pe99_35(.x(x35),.w(w99_34),.acc(r99_34),.res(r99_35),.clk(clk),.wout(w99_35));
	PE pe99_36(.x(x36),.w(w99_35),.acc(r99_35),.res(r99_36),.clk(clk),.wout(w99_36));
	PE pe99_37(.x(x37),.w(w99_36),.acc(r99_36),.res(r99_37),.clk(clk),.wout(w99_37));
	PE pe99_38(.x(x38),.w(w99_37),.acc(r99_37),.res(r99_38),.clk(clk),.wout(w99_38));
	PE pe99_39(.x(x39),.w(w99_38),.acc(r99_38),.res(r99_39),.clk(clk),.wout(w99_39));
	PE pe99_40(.x(x40),.w(w99_39),.acc(r99_39),.res(r99_40),.clk(clk),.wout(w99_40));
	PE pe99_41(.x(x41),.w(w99_40),.acc(r99_40),.res(r99_41),.clk(clk),.wout(w99_41));
	PE pe99_42(.x(x42),.w(w99_41),.acc(r99_41),.res(r99_42),.clk(clk),.wout(w99_42));
	PE pe99_43(.x(x43),.w(w99_42),.acc(r99_42),.res(r99_43),.clk(clk),.wout(w99_43));
	PE pe99_44(.x(x44),.w(w99_43),.acc(r99_43),.res(r99_44),.clk(clk),.wout(w99_44));
	PE pe99_45(.x(x45),.w(w99_44),.acc(r99_44),.res(r99_45),.clk(clk),.wout(w99_45));
	PE pe99_46(.x(x46),.w(w99_45),.acc(r99_45),.res(r99_46),.clk(clk),.wout(w99_46));
	PE pe99_47(.x(x47),.w(w99_46),.acc(r99_46),.res(r99_47),.clk(clk),.wout(w99_47));
	PE pe99_48(.x(x48),.w(w99_47),.acc(r99_47),.res(r99_48),.clk(clk),.wout(w99_48));
	PE pe99_49(.x(x49),.w(w99_48),.acc(r99_48),.res(r99_49),.clk(clk),.wout(w99_49));
	PE pe99_50(.x(x50),.w(w99_49),.acc(r99_49),.res(r99_50),.clk(clk),.wout(w99_50));
	PE pe99_51(.x(x51),.w(w99_50),.acc(r99_50),.res(r99_51),.clk(clk),.wout(w99_51));
	PE pe99_52(.x(x52),.w(w99_51),.acc(r99_51),.res(r99_52),.clk(clk),.wout(w99_52));
	PE pe99_53(.x(x53),.w(w99_52),.acc(r99_52),.res(r99_53),.clk(clk),.wout(w99_53));
	PE pe99_54(.x(x54),.w(w99_53),.acc(r99_53),.res(r99_54),.clk(clk),.wout(w99_54));
	PE pe99_55(.x(x55),.w(w99_54),.acc(r99_54),.res(r99_55),.clk(clk),.wout(w99_55));
	PE pe99_56(.x(x56),.w(w99_55),.acc(r99_55),.res(r99_56),.clk(clk),.wout(w99_56));
	PE pe99_57(.x(x57),.w(w99_56),.acc(r99_56),.res(r99_57),.clk(clk),.wout(w99_57));
	PE pe99_58(.x(x58),.w(w99_57),.acc(r99_57),.res(r99_58),.clk(clk),.wout(w99_58));
	PE pe99_59(.x(x59),.w(w99_58),.acc(r99_58),.res(r99_59),.clk(clk),.wout(w99_59));
	PE pe99_60(.x(x60),.w(w99_59),.acc(r99_59),.res(r99_60),.clk(clk),.wout(w99_60));
	PE pe99_61(.x(x61),.w(w99_60),.acc(r99_60),.res(r99_61),.clk(clk),.wout(w99_61));
	PE pe99_62(.x(x62),.w(w99_61),.acc(r99_61),.res(r99_62),.clk(clk),.wout(w99_62));
	PE pe99_63(.x(x63),.w(w99_62),.acc(r99_62),.res(r99_63),.clk(clk),.wout(w99_63));
	PE pe99_64(.x(x64),.w(w99_63),.acc(r99_63),.res(r99_64),.clk(clk),.wout(w99_64));
	PE pe99_65(.x(x65),.w(w99_64),.acc(r99_64),.res(r99_65),.clk(clk),.wout(w99_65));
	PE pe99_66(.x(x66),.w(w99_65),.acc(r99_65),.res(r99_66),.clk(clk),.wout(w99_66));
	PE pe99_67(.x(x67),.w(w99_66),.acc(r99_66),.res(r99_67),.clk(clk),.wout(w99_67));
	PE pe99_68(.x(x68),.w(w99_67),.acc(r99_67),.res(r99_68),.clk(clk),.wout(w99_68));
	PE pe99_69(.x(x69),.w(w99_68),.acc(r99_68),.res(r99_69),.clk(clk),.wout(w99_69));
	PE pe99_70(.x(x70),.w(w99_69),.acc(r99_69),.res(r99_70),.clk(clk),.wout(w99_70));
	PE pe99_71(.x(x71),.w(w99_70),.acc(r99_70),.res(r99_71),.clk(clk),.wout(w99_71));
	PE pe99_72(.x(x72),.w(w99_71),.acc(r99_71),.res(r99_72),.clk(clk),.wout(w99_72));
	PE pe99_73(.x(x73),.w(w99_72),.acc(r99_72),.res(r99_73),.clk(clk),.wout(w99_73));
	PE pe99_74(.x(x74),.w(w99_73),.acc(r99_73),.res(r99_74),.clk(clk),.wout(w99_74));
	PE pe99_75(.x(x75),.w(w99_74),.acc(r99_74),.res(r99_75),.clk(clk),.wout(w99_75));
	PE pe99_76(.x(x76),.w(w99_75),.acc(r99_75),.res(r99_76),.clk(clk),.wout(w99_76));
	PE pe99_77(.x(x77),.w(w99_76),.acc(r99_76),.res(r99_77),.clk(clk),.wout(w99_77));
	PE pe99_78(.x(x78),.w(w99_77),.acc(r99_77),.res(r99_78),.clk(clk),.wout(w99_78));
	PE pe99_79(.x(x79),.w(w99_78),.acc(r99_78),.res(r99_79),.clk(clk),.wout(w99_79));
	PE pe99_80(.x(x80),.w(w99_79),.acc(r99_79),.res(r99_80),.clk(clk),.wout(w99_80));
	PE pe99_81(.x(x81),.w(w99_80),.acc(r99_80),.res(r99_81),.clk(clk),.wout(w99_81));
	PE pe99_82(.x(x82),.w(w99_81),.acc(r99_81),.res(r99_82),.clk(clk),.wout(w99_82));
	PE pe99_83(.x(x83),.w(w99_82),.acc(r99_82),.res(r99_83),.clk(clk),.wout(w99_83));
	PE pe99_84(.x(x84),.w(w99_83),.acc(r99_83),.res(r99_84),.clk(clk),.wout(w99_84));
	PE pe99_85(.x(x85),.w(w99_84),.acc(r99_84),.res(r99_85),.clk(clk),.wout(w99_85));
	PE pe99_86(.x(x86),.w(w99_85),.acc(r99_85),.res(r99_86),.clk(clk),.wout(w99_86));
	PE pe99_87(.x(x87),.w(w99_86),.acc(r99_86),.res(r99_87),.clk(clk),.wout(w99_87));
	PE pe99_88(.x(x88),.w(w99_87),.acc(r99_87),.res(r99_88),.clk(clk),.wout(w99_88));
	PE pe99_89(.x(x89),.w(w99_88),.acc(r99_88),.res(r99_89),.clk(clk),.wout(w99_89));
	PE pe99_90(.x(x90),.w(w99_89),.acc(r99_89),.res(r99_90),.clk(clk),.wout(w99_90));
	PE pe99_91(.x(x91),.w(w99_90),.acc(r99_90),.res(r99_91),.clk(clk),.wout(w99_91));
	PE pe99_92(.x(x92),.w(w99_91),.acc(r99_91),.res(r99_92),.clk(clk),.wout(w99_92));
	PE pe99_93(.x(x93),.w(w99_92),.acc(r99_92),.res(r99_93),.clk(clk),.wout(w99_93));
	PE pe99_94(.x(x94),.w(w99_93),.acc(r99_93),.res(r99_94),.clk(clk),.wout(w99_94));
	PE pe99_95(.x(x95),.w(w99_94),.acc(r99_94),.res(r99_95),.clk(clk),.wout(w99_95));
	PE pe99_96(.x(x96),.w(w99_95),.acc(r99_95),.res(r99_96),.clk(clk),.wout(w99_96));
	PE pe99_97(.x(x97),.w(w99_96),.acc(r99_96),.res(r99_97),.clk(clk),.wout(w99_97));
	PE pe99_98(.x(x98),.w(w99_97),.acc(r99_97),.res(r99_98),.clk(clk),.wout(w99_98));
	PE pe99_99(.x(x99),.w(w99_98),.acc(r99_98),.res(r99_99),.clk(clk),.wout(w99_99));
	PE pe99_100(.x(x100),.w(w99_99),.acc(r99_99),.res(r99_100),.clk(clk),.wout(w99_100));
	PE pe99_101(.x(x101),.w(w99_100),.acc(r99_100),.res(r99_101),.clk(clk),.wout(w99_101));
	PE pe99_102(.x(x102),.w(w99_101),.acc(r99_101),.res(r99_102),.clk(clk),.wout(w99_102));
	PE pe99_103(.x(x103),.w(w99_102),.acc(r99_102),.res(r99_103),.clk(clk),.wout(w99_103));
	PE pe99_104(.x(x104),.w(w99_103),.acc(r99_103),.res(r99_104),.clk(clk),.wout(w99_104));
	PE pe99_105(.x(x105),.w(w99_104),.acc(r99_104),.res(r99_105),.clk(clk),.wout(w99_105));
	PE pe99_106(.x(x106),.w(w99_105),.acc(r99_105),.res(r99_106),.clk(clk),.wout(w99_106));
	PE pe99_107(.x(x107),.w(w99_106),.acc(r99_106),.res(r99_107),.clk(clk),.wout(w99_107));
	PE pe99_108(.x(x108),.w(w99_107),.acc(r99_107),.res(r99_108),.clk(clk),.wout(w99_108));
	PE pe99_109(.x(x109),.w(w99_108),.acc(r99_108),.res(r99_109),.clk(clk),.wout(w99_109));
	PE pe99_110(.x(x110),.w(w99_109),.acc(r99_109),.res(r99_110),.clk(clk),.wout(w99_110));
	PE pe99_111(.x(x111),.w(w99_110),.acc(r99_110),.res(r99_111),.clk(clk),.wout(w99_111));
	PE pe99_112(.x(x112),.w(w99_111),.acc(r99_111),.res(r99_112),.clk(clk),.wout(w99_112));
	PE pe99_113(.x(x113),.w(w99_112),.acc(r99_112),.res(r99_113),.clk(clk),.wout(w99_113));
	PE pe99_114(.x(x114),.w(w99_113),.acc(r99_113),.res(r99_114),.clk(clk),.wout(w99_114));
	PE pe99_115(.x(x115),.w(w99_114),.acc(r99_114),.res(r99_115),.clk(clk),.wout(w99_115));
	PE pe99_116(.x(x116),.w(w99_115),.acc(r99_115),.res(r99_116),.clk(clk),.wout(w99_116));
	PE pe99_117(.x(x117),.w(w99_116),.acc(r99_116),.res(r99_117),.clk(clk),.wout(w99_117));
	PE pe99_118(.x(x118),.w(w99_117),.acc(r99_117),.res(r99_118),.clk(clk),.wout(w99_118));
	PE pe99_119(.x(x119),.w(w99_118),.acc(r99_118),.res(r99_119),.clk(clk),.wout(w99_119));
	PE pe99_120(.x(x120),.w(w99_119),.acc(r99_119),.res(r99_120),.clk(clk),.wout(w99_120));
	PE pe99_121(.x(x121),.w(w99_120),.acc(r99_120),.res(r99_121),.clk(clk),.wout(w99_121));
	PE pe99_122(.x(x122),.w(w99_121),.acc(r99_121),.res(r99_122),.clk(clk),.wout(w99_122));
	PE pe99_123(.x(x123),.w(w99_122),.acc(r99_122),.res(r99_123),.clk(clk),.wout(w99_123));
	PE pe99_124(.x(x124),.w(w99_123),.acc(r99_123),.res(r99_124),.clk(clk),.wout(w99_124));
	PE pe99_125(.x(x125),.w(w99_124),.acc(r99_124),.res(r99_125),.clk(clk),.wout(w99_125));
	PE pe99_126(.x(x126),.w(w99_125),.acc(r99_125),.res(r99_126),.clk(clk),.wout(w99_126));
	PE pe99_127(.x(x127),.w(w99_126),.acc(r99_126),.res(result99),.clk(clk),.wout(weight99));

	PE pe100_0(.x(x0),.w(w100),.acc(32'h0),.res(r100_0),.clk(clk),.wout(w100_0));
	PE pe100_1(.x(x1),.w(w100_0),.acc(r100_0),.res(r100_1),.clk(clk),.wout(w100_1));
	PE pe100_2(.x(x2),.w(w100_1),.acc(r100_1),.res(r100_2),.clk(clk),.wout(w100_2));
	PE pe100_3(.x(x3),.w(w100_2),.acc(r100_2),.res(r100_3),.clk(clk),.wout(w100_3));
	PE pe100_4(.x(x4),.w(w100_3),.acc(r100_3),.res(r100_4),.clk(clk),.wout(w100_4));
	PE pe100_5(.x(x5),.w(w100_4),.acc(r100_4),.res(r100_5),.clk(clk),.wout(w100_5));
	PE pe100_6(.x(x6),.w(w100_5),.acc(r100_5),.res(r100_6),.clk(clk),.wout(w100_6));
	PE pe100_7(.x(x7),.w(w100_6),.acc(r100_6),.res(r100_7),.clk(clk),.wout(w100_7));
	PE pe100_8(.x(x8),.w(w100_7),.acc(r100_7),.res(r100_8),.clk(clk),.wout(w100_8));
	PE pe100_9(.x(x9),.w(w100_8),.acc(r100_8),.res(r100_9),.clk(clk),.wout(w100_9));
	PE pe100_10(.x(x10),.w(w100_9),.acc(r100_9),.res(r100_10),.clk(clk),.wout(w100_10));
	PE pe100_11(.x(x11),.w(w100_10),.acc(r100_10),.res(r100_11),.clk(clk),.wout(w100_11));
	PE pe100_12(.x(x12),.w(w100_11),.acc(r100_11),.res(r100_12),.clk(clk),.wout(w100_12));
	PE pe100_13(.x(x13),.w(w100_12),.acc(r100_12),.res(r100_13),.clk(clk),.wout(w100_13));
	PE pe100_14(.x(x14),.w(w100_13),.acc(r100_13),.res(r100_14),.clk(clk),.wout(w100_14));
	PE pe100_15(.x(x15),.w(w100_14),.acc(r100_14),.res(r100_15),.clk(clk),.wout(w100_15));
	PE pe100_16(.x(x16),.w(w100_15),.acc(r100_15),.res(r100_16),.clk(clk),.wout(w100_16));
	PE pe100_17(.x(x17),.w(w100_16),.acc(r100_16),.res(r100_17),.clk(clk),.wout(w100_17));
	PE pe100_18(.x(x18),.w(w100_17),.acc(r100_17),.res(r100_18),.clk(clk),.wout(w100_18));
	PE pe100_19(.x(x19),.w(w100_18),.acc(r100_18),.res(r100_19),.clk(clk),.wout(w100_19));
	PE pe100_20(.x(x20),.w(w100_19),.acc(r100_19),.res(r100_20),.clk(clk),.wout(w100_20));
	PE pe100_21(.x(x21),.w(w100_20),.acc(r100_20),.res(r100_21),.clk(clk),.wout(w100_21));
	PE pe100_22(.x(x22),.w(w100_21),.acc(r100_21),.res(r100_22),.clk(clk),.wout(w100_22));
	PE pe100_23(.x(x23),.w(w100_22),.acc(r100_22),.res(r100_23),.clk(clk),.wout(w100_23));
	PE pe100_24(.x(x24),.w(w100_23),.acc(r100_23),.res(r100_24),.clk(clk),.wout(w100_24));
	PE pe100_25(.x(x25),.w(w100_24),.acc(r100_24),.res(r100_25),.clk(clk),.wout(w100_25));
	PE pe100_26(.x(x26),.w(w100_25),.acc(r100_25),.res(r100_26),.clk(clk),.wout(w100_26));
	PE pe100_27(.x(x27),.w(w100_26),.acc(r100_26),.res(r100_27),.clk(clk),.wout(w100_27));
	PE pe100_28(.x(x28),.w(w100_27),.acc(r100_27),.res(r100_28),.clk(clk),.wout(w100_28));
	PE pe100_29(.x(x29),.w(w100_28),.acc(r100_28),.res(r100_29),.clk(clk),.wout(w100_29));
	PE pe100_30(.x(x30),.w(w100_29),.acc(r100_29),.res(r100_30),.clk(clk),.wout(w100_30));
	PE pe100_31(.x(x31),.w(w100_30),.acc(r100_30),.res(r100_31),.clk(clk),.wout(w100_31));
	PE pe100_32(.x(x32),.w(w100_31),.acc(r100_31),.res(r100_32),.clk(clk),.wout(w100_32));
	PE pe100_33(.x(x33),.w(w100_32),.acc(r100_32),.res(r100_33),.clk(clk),.wout(w100_33));
	PE pe100_34(.x(x34),.w(w100_33),.acc(r100_33),.res(r100_34),.clk(clk),.wout(w100_34));
	PE pe100_35(.x(x35),.w(w100_34),.acc(r100_34),.res(r100_35),.clk(clk),.wout(w100_35));
	PE pe100_36(.x(x36),.w(w100_35),.acc(r100_35),.res(r100_36),.clk(clk),.wout(w100_36));
	PE pe100_37(.x(x37),.w(w100_36),.acc(r100_36),.res(r100_37),.clk(clk),.wout(w100_37));
	PE pe100_38(.x(x38),.w(w100_37),.acc(r100_37),.res(r100_38),.clk(clk),.wout(w100_38));
	PE pe100_39(.x(x39),.w(w100_38),.acc(r100_38),.res(r100_39),.clk(clk),.wout(w100_39));
	PE pe100_40(.x(x40),.w(w100_39),.acc(r100_39),.res(r100_40),.clk(clk),.wout(w100_40));
	PE pe100_41(.x(x41),.w(w100_40),.acc(r100_40),.res(r100_41),.clk(clk),.wout(w100_41));
	PE pe100_42(.x(x42),.w(w100_41),.acc(r100_41),.res(r100_42),.clk(clk),.wout(w100_42));
	PE pe100_43(.x(x43),.w(w100_42),.acc(r100_42),.res(r100_43),.clk(clk),.wout(w100_43));
	PE pe100_44(.x(x44),.w(w100_43),.acc(r100_43),.res(r100_44),.clk(clk),.wout(w100_44));
	PE pe100_45(.x(x45),.w(w100_44),.acc(r100_44),.res(r100_45),.clk(clk),.wout(w100_45));
	PE pe100_46(.x(x46),.w(w100_45),.acc(r100_45),.res(r100_46),.clk(clk),.wout(w100_46));
	PE pe100_47(.x(x47),.w(w100_46),.acc(r100_46),.res(r100_47),.clk(clk),.wout(w100_47));
	PE pe100_48(.x(x48),.w(w100_47),.acc(r100_47),.res(r100_48),.clk(clk),.wout(w100_48));
	PE pe100_49(.x(x49),.w(w100_48),.acc(r100_48),.res(r100_49),.clk(clk),.wout(w100_49));
	PE pe100_50(.x(x50),.w(w100_49),.acc(r100_49),.res(r100_50),.clk(clk),.wout(w100_50));
	PE pe100_51(.x(x51),.w(w100_50),.acc(r100_50),.res(r100_51),.clk(clk),.wout(w100_51));
	PE pe100_52(.x(x52),.w(w100_51),.acc(r100_51),.res(r100_52),.clk(clk),.wout(w100_52));
	PE pe100_53(.x(x53),.w(w100_52),.acc(r100_52),.res(r100_53),.clk(clk),.wout(w100_53));
	PE pe100_54(.x(x54),.w(w100_53),.acc(r100_53),.res(r100_54),.clk(clk),.wout(w100_54));
	PE pe100_55(.x(x55),.w(w100_54),.acc(r100_54),.res(r100_55),.clk(clk),.wout(w100_55));
	PE pe100_56(.x(x56),.w(w100_55),.acc(r100_55),.res(r100_56),.clk(clk),.wout(w100_56));
	PE pe100_57(.x(x57),.w(w100_56),.acc(r100_56),.res(r100_57),.clk(clk),.wout(w100_57));
	PE pe100_58(.x(x58),.w(w100_57),.acc(r100_57),.res(r100_58),.clk(clk),.wout(w100_58));
	PE pe100_59(.x(x59),.w(w100_58),.acc(r100_58),.res(r100_59),.clk(clk),.wout(w100_59));
	PE pe100_60(.x(x60),.w(w100_59),.acc(r100_59),.res(r100_60),.clk(clk),.wout(w100_60));
	PE pe100_61(.x(x61),.w(w100_60),.acc(r100_60),.res(r100_61),.clk(clk),.wout(w100_61));
	PE pe100_62(.x(x62),.w(w100_61),.acc(r100_61),.res(r100_62),.clk(clk),.wout(w100_62));
	PE pe100_63(.x(x63),.w(w100_62),.acc(r100_62),.res(r100_63),.clk(clk),.wout(w100_63));
	PE pe100_64(.x(x64),.w(w100_63),.acc(r100_63),.res(r100_64),.clk(clk),.wout(w100_64));
	PE pe100_65(.x(x65),.w(w100_64),.acc(r100_64),.res(r100_65),.clk(clk),.wout(w100_65));
	PE pe100_66(.x(x66),.w(w100_65),.acc(r100_65),.res(r100_66),.clk(clk),.wout(w100_66));
	PE pe100_67(.x(x67),.w(w100_66),.acc(r100_66),.res(r100_67),.clk(clk),.wout(w100_67));
	PE pe100_68(.x(x68),.w(w100_67),.acc(r100_67),.res(r100_68),.clk(clk),.wout(w100_68));
	PE pe100_69(.x(x69),.w(w100_68),.acc(r100_68),.res(r100_69),.clk(clk),.wout(w100_69));
	PE pe100_70(.x(x70),.w(w100_69),.acc(r100_69),.res(r100_70),.clk(clk),.wout(w100_70));
	PE pe100_71(.x(x71),.w(w100_70),.acc(r100_70),.res(r100_71),.clk(clk),.wout(w100_71));
	PE pe100_72(.x(x72),.w(w100_71),.acc(r100_71),.res(r100_72),.clk(clk),.wout(w100_72));
	PE pe100_73(.x(x73),.w(w100_72),.acc(r100_72),.res(r100_73),.clk(clk),.wout(w100_73));
	PE pe100_74(.x(x74),.w(w100_73),.acc(r100_73),.res(r100_74),.clk(clk),.wout(w100_74));
	PE pe100_75(.x(x75),.w(w100_74),.acc(r100_74),.res(r100_75),.clk(clk),.wout(w100_75));
	PE pe100_76(.x(x76),.w(w100_75),.acc(r100_75),.res(r100_76),.clk(clk),.wout(w100_76));
	PE pe100_77(.x(x77),.w(w100_76),.acc(r100_76),.res(r100_77),.clk(clk),.wout(w100_77));
	PE pe100_78(.x(x78),.w(w100_77),.acc(r100_77),.res(r100_78),.clk(clk),.wout(w100_78));
	PE pe100_79(.x(x79),.w(w100_78),.acc(r100_78),.res(r100_79),.clk(clk),.wout(w100_79));
	PE pe100_80(.x(x80),.w(w100_79),.acc(r100_79),.res(r100_80),.clk(clk),.wout(w100_80));
	PE pe100_81(.x(x81),.w(w100_80),.acc(r100_80),.res(r100_81),.clk(clk),.wout(w100_81));
	PE pe100_82(.x(x82),.w(w100_81),.acc(r100_81),.res(r100_82),.clk(clk),.wout(w100_82));
	PE pe100_83(.x(x83),.w(w100_82),.acc(r100_82),.res(r100_83),.clk(clk),.wout(w100_83));
	PE pe100_84(.x(x84),.w(w100_83),.acc(r100_83),.res(r100_84),.clk(clk),.wout(w100_84));
	PE pe100_85(.x(x85),.w(w100_84),.acc(r100_84),.res(r100_85),.clk(clk),.wout(w100_85));
	PE pe100_86(.x(x86),.w(w100_85),.acc(r100_85),.res(r100_86),.clk(clk),.wout(w100_86));
	PE pe100_87(.x(x87),.w(w100_86),.acc(r100_86),.res(r100_87),.clk(clk),.wout(w100_87));
	PE pe100_88(.x(x88),.w(w100_87),.acc(r100_87),.res(r100_88),.clk(clk),.wout(w100_88));
	PE pe100_89(.x(x89),.w(w100_88),.acc(r100_88),.res(r100_89),.clk(clk),.wout(w100_89));
	PE pe100_90(.x(x90),.w(w100_89),.acc(r100_89),.res(r100_90),.clk(clk),.wout(w100_90));
	PE pe100_91(.x(x91),.w(w100_90),.acc(r100_90),.res(r100_91),.clk(clk),.wout(w100_91));
	PE pe100_92(.x(x92),.w(w100_91),.acc(r100_91),.res(r100_92),.clk(clk),.wout(w100_92));
	PE pe100_93(.x(x93),.w(w100_92),.acc(r100_92),.res(r100_93),.clk(clk),.wout(w100_93));
	PE pe100_94(.x(x94),.w(w100_93),.acc(r100_93),.res(r100_94),.clk(clk),.wout(w100_94));
	PE pe100_95(.x(x95),.w(w100_94),.acc(r100_94),.res(r100_95),.clk(clk),.wout(w100_95));
	PE pe100_96(.x(x96),.w(w100_95),.acc(r100_95),.res(r100_96),.clk(clk),.wout(w100_96));
	PE pe100_97(.x(x97),.w(w100_96),.acc(r100_96),.res(r100_97),.clk(clk),.wout(w100_97));
	PE pe100_98(.x(x98),.w(w100_97),.acc(r100_97),.res(r100_98),.clk(clk),.wout(w100_98));
	PE pe100_99(.x(x99),.w(w100_98),.acc(r100_98),.res(r100_99),.clk(clk),.wout(w100_99));
	PE pe100_100(.x(x100),.w(w100_99),.acc(r100_99),.res(r100_100),.clk(clk),.wout(w100_100));
	PE pe100_101(.x(x101),.w(w100_100),.acc(r100_100),.res(r100_101),.clk(clk),.wout(w100_101));
	PE pe100_102(.x(x102),.w(w100_101),.acc(r100_101),.res(r100_102),.clk(clk),.wout(w100_102));
	PE pe100_103(.x(x103),.w(w100_102),.acc(r100_102),.res(r100_103),.clk(clk),.wout(w100_103));
	PE pe100_104(.x(x104),.w(w100_103),.acc(r100_103),.res(r100_104),.clk(clk),.wout(w100_104));
	PE pe100_105(.x(x105),.w(w100_104),.acc(r100_104),.res(r100_105),.clk(clk),.wout(w100_105));
	PE pe100_106(.x(x106),.w(w100_105),.acc(r100_105),.res(r100_106),.clk(clk),.wout(w100_106));
	PE pe100_107(.x(x107),.w(w100_106),.acc(r100_106),.res(r100_107),.clk(clk),.wout(w100_107));
	PE pe100_108(.x(x108),.w(w100_107),.acc(r100_107),.res(r100_108),.clk(clk),.wout(w100_108));
	PE pe100_109(.x(x109),.w(w100_108),.acc(r100_108),.res(r100_109),.clk(clk),.wout(w100_109));
	PE pe100_110(.x(x110),.w(w100_109),.acc(r100_109),.res(r100_110),.clk(clk),.wout(w100_110));
	PE pe100_111(.x(x111),.w(w100_110),.acc(r100_110),.res(r100_111),.clk(clk),.wout(w100_111));
	PE pe100_112(.x(x112),.w(w100_111),.acc(r100_111),.res(r100_112),.clk(clk),.wout(w100_112));
	PE pe100_113(.x(x113),.w(w100_112),.acc(r100_112),.res(r100_113),.clk(clk),.wout(w100_113));
	PE pe100_114(.x(x114),.w(w100_113),.acc(r100_113),.res(r100_114),.clk(clk),.wout(w100_114));
	PE pe100_115(.x(x115),.w(w100_114),.acc(r100_114),.res(r100_115),.clk(clk),.wout(w100_115));
	PE pe100_116(.x(x116),.w(w100_115),.acc(r100_115),.res(r100_116),.clk(clk),.wout(w100_116));
	PE pe100_117(.x(x117),.w(w100_116),.acc(r100_116),.res(r100_117),.clk(clk),.wout(w100_117));
	PE pe100_118(.x(x118),.w(w100_117),.acc(r100_117),.res(r100_118),.clk(clk),.wout(w100_118));
	PE pe100_119(.x(x119),.w(w100_118),.acc(r100_118),.res(r100_119),.clk(clk),.wout(w100_119));
	PE pe100_120(.x(x120),.w(w100_119),.acc(r100_119),.res(r100_120),.clk(clk),.wout(w100_120));
	PE pe100_121(.x(x121),.w(w100_120),.acc(r100_120),.res(r100_121),.clk(clk),.wout(w100_121));
	PE pe100_122(.x(x122),.w(w100_121),.acc(r100_121),.res(r100_122),.clk(clk),.wout(w100_122));
	PE pe100_123(.x(x123),.w(w100_122),.acc(r100_122),.res(r100_123),.clk(clk),.wout(w100_123));
	PE pe100_124(.x(x124),.w(w100_123),.acc(r100_123),.res(r100_124),.clk(clk),.wout(w100_124));
	PE pe100_125(.x(x125),.w(w100_124),.acc(r100_124),.res(r100_125),.clk(clk),.wout(w100_125));
	PE pe100_126(.x(x126),.w(w100_125),.acc(r100_125),.res(r100_126),.clk(clk),.wout(w100_126));
	PE pe100_127(.x(x127),.w(w100_126),.acc(r100_126),.res(result100),.clk(clk),.wout(weight100));

	PE pe101_0(.x(x0),.w(w101),.acc(32'h0),.res(r101_0),.clk(clk),.wout(w101_0));
	PE pe101_1(.x(x1),.w(w101_0),.acc(r101_0),.res(r101_1),.clk(clk),.wout(w101_1));
	PE pe101_2(.x(x2),.w(w101_1),.acc(r101_1),.res(r101_2),.clk(clk),.wout(w101_2));
	PE pe101_3(.x(x3),.w(w101_2),.acc(r101_2),.res(r101_3),.clk(clk),.wout(w101_3));
	PE pe101_4(.x(x4),.w(w101_3),.acc(r101_3),.res(r101_4),.clk(clk),.wout(w101_4));
	PE pe101_5(.x(x5),.w(w101_4),.acc(r101_4),.res(r101_5),.clk(clk),.wout(w101_5));
	PE pe101_6(.x(x6),.w(w101_5),.acc(r101_5),.res(r101_6),.clk(clk),.wout(w101_6));
	PE pe101_7(.x(x7),.w(w101_6),.acc(r101_6),.res(r101_7),.clk(clk),.wout(w101_7));
	PE pe101_8(.x(x8),.w(w101_7),.acc(r101_7),.res(r101_8),.clk(clk),.wout(w101_8));
	PE pe101_9(.x(x9),.w(w101_8),.acc(r101_8),.res(r101_9),.clk(clk),.wout(w101_9));
	PE pe101_10(.x(x10),.w(w101_9),.acc(r101_9),.res(r101_10),.clk(clk),.wout(w101_10));
	PE pe101_11(.x(x11),.w(w101_10),.acc(r101_10),.res(r101_11),.clk(clk),.wout(w101_11));
	PE pe101_12(.x(x12),.w(w101_11),.acc(r101_11),.res(r101_12),.clk(clk),.wout(w101_12));
	PE pe101_13(.x(x13),.w(w101_12),.acc(r101_12),.res(r101_13),.clk(clk),.wout(w101_13));
	PE pe101_14(.x(x14),.w(w101_13),.acc(r101_13),.res(r101_14),.clk(clk),.wout(w101_14));
	PE pe101_15(.x(x15),.w(w101_14),.acc(r101_14),.res(r101_15),.clk(clk),.wout(w101_15));
	PE pe101_16(.x(x16),.w(w101_15),.acc(r101_15),.res(r101_16),.clk(clk),.wout(w101_16));
	PE pe101_17(.x(x17),.w(w101_16),.acc(r101_16),.res(r101_17),.clk(clk),.wout(w101_17));
	PE pe101_18(.x(x18),.w(w101_17),.acc(r101_17),.res(r101_18),.clk(clk),.wout(w101_18));
	PE pe101_19(.x(x19),.w(w101_18),.acc(r101_18),.res(r101_19),.clk(clk),.wout(w101_19));
	PE pe101_20(.x(x20),.w(w101_19),.acc(r101_19),.res(r101_20),.clk(clk),.wout(w101_20));
	PE pe101_21(.x(x21),.w(w101_20),.acc(r101_20),.res(r101_21),.clk(clk),.wout(w101_21));
	PE pe101_22(.x(x22),.w(w101_21),.acc(r101_21),.res(r101_22),.clk(clk),.wout(w101_22));
	PE pe101_23(.x(x23),.w(w101_22),.acc(r101_22),.res(r101_23),.clk(clk),.wout(w101_23));
	PE pe101_24(.x(x24),.w(w101_23),.acc(r101_23),.res(r101_24),.clk(clk),.wout(w101_24));
	PE pe101_25(.x(x25),.w(w101_24),.acc(r101_24),.res(r101_25),.clk(clk),.wout(w101_25));
	PE pe101_26(.x(x26),.w(w101_25),.acc(r101_25),.res(r101_26),.clk(clk),.wout(w101_26));
	PE pe101_27(.x(x27),.w(w101_26),.acc(r101_26),.res(r101_27),.clk(clk),.wout(w101_27));
	PE pe101_28(.x(x28),.w(w101_27),.acc(r101_27),.res(r101_28),.clk(clk),.wout(w101_28));
	PE pe101_29(.x(x29),.w(w101_28),.acc(r101_28),.res(r101_29),.clk(clk),.wout(w101_29));
	PE pe101_30(.x(x30),.w(w101_29),.acc(r101_29),.res(r101_30),.clk(clk),.wout(w101_30));
	PE pe101_31(.x(x31),.w(w101_30),.acc(r101_30),.res(r101_31),.clk(clk),.wout(w101_31));
	PE pe101_32(.x(x32),.w(w101_31),.acc(r101_31),.res(r101_32),.clk(clk),.wout(w101_32));
	PE pe101_33(.x(x33),.w(w101_32),.acc(r101_32),.res(r101_33),.clk(clk),.wout(w101_33));
	PE pe101_34(.x(x34),.w(w101_33),.acc(r101_33),.res(r101_34),.clk(clk),.wout(w101_34));
	PE pe101_35(.x(x35),.w(w101_34),.acc(r101_34),.res(r101_35),.clk(clk),.wout(w101_35));
	PE pe101_36(.x(x36),.w(w101_35),.acc(r101_35),.res(r101_36),.clk(clk),.wout(w101_36));
	PE pe101_37(.x(x37),.w(w101_36),.acc(r101_36),.res(r101_37),.clk(clk),.wout(w101_37));
	PE pe101_38(.x(x38),.w(w101_37),.acc(r101_37),.res(r101_38),.clk(clk),.wout(w101_38));
	PE pe101_39(.x(x39),.w(w101_38),.acc(r101_38),.res(r101_39),.clk(clk),.wout(w101_39));
	PE pe101_40(.x(x40),.w(w101_39),.acc(r101_39),.res(r101_40),.clk(clk),.wout(w101_40));
	PE pe101_41(.x(x41),.w(w101_40),.acc(r101_40),.res(r101_41),.clk(clk),.wout(w101_41));
	PE pe101_42(.x(x42),.w(w101_41),.acc(r101_41),.res(r101_42),.clk(clk),.wout(w101_42));
	PE pe101_43(.x(x43),.w(w101_42),.acc(r101_42),.res(r101_43),.clk(clk),.wout(w101_43));
	PE pe101_44(.x(x44),.w(w101_43),.acc(r101_43),.res(r101_44),.clk(clk),.wout(w101_44));
	PE pe101_45(.x(x45),.w(w101_44),.acc(r101_44),.res(r101_45),.clk(clk),.wout(w101_45));
	PE pe101_46(.x(x46),.w(w101_45),.acc(r101_45),.res(r101_46),.clk(clk),.wout(w101_46));
	PE pe101_47(.x(x47),.w(w101_46),.acc(r101_46),.res(r101_47),.clk(clk),.wout(w101_47));
	PE pe101_48(.x(x48),.w(w101_47),.acc(r101_47),.res(r101_48),.clk(clk),.wout(w101_48));
	PE pe101_49(.x(x49),.w(w101_48),.acc(r101_48),.res(r101_49),.clk(clk),.wout(w101_49));
	PE pe101_50(.x(x50),.w(w101_49),.acc(r101_49),.res(r101_50),.clk(clk),.wout(w101_50));
	PE pe101_51(.x(x51),.w(w101_50),.acc(r101_50),.res(r101_51),.clk(clk),.wout(w101_51));
	PE pe101_52(.x(x52),.w(w101_51),.acc(r101_51),.res(r101_52),.clk(clk),.wout(w101_52));
	PE pe101_53(.x(x53),.w(w101_52),.acc(r101_52),.res(r101_53),.clk(clk),.wout(w101_53));
	PE pe101_54(.x(x54),.w(w101_53),.acc(r101_53),.res(r101_54),.clk(clk),.wout(w101_54));
	PE pe101_55(.x(x55),.w(w101_54),.acc(r101_54),.res(r101_55),.clk(clk),.wout(w101_55));
	PE pe101_56(.x(x56),.w(w101_55),.acc(r101_55),.res(r101_56),.clk(clk),.wout(w101_56));
	PE pe101_57(.x(x57),.w(w101_56),.acc(r101_56),.res(r101_57),.clk(clk),.wout(w101_57));
	PE pe101_58(.x(x58),.w(w101_57),.acc(r101_57),.res(r101_58),.clk(clk),.wout(w101_58));
	PE pe101_59(.x(x59),.w(w101_58),.acc(r101_58),.res(r101_59),.clk(clk),.wout(w101_59));
	PE pe101_60(.x(x60),.w(w101_59),.acc(r101_59),.res(r101_60),.clk(clk),.wout(w101_60));
	PE pe101_61(.x(x61),.w(w101_60),.acc(r101_60),.res(r101_61),.clk(clk),.wout(w101_61));
	PE pe101_62(.x(x62),.w(w101_61),.acc(r101_61),.res(r101_62),.clk(clk),.wout(w101_62));
	PE pe101_63(.x(x63),.w(w101_62),.acc(r101_62),.res(r101_63),.clk(clk),.wout(w101_63));
	PE pe101_64(.x(x64),.w(w101_63),.acc(r101_63),.res(r101_64),.clk(clk),.wout(w101_64));
	PE pe101_65(.x(x65),.w(w101_64),.acc(r101_64),.res(r101_65),.clk(clk),.wout(w101_65));
	PE pe101_66(.x(x66),.w(w101_65),.acc(r101_65),.res(r101_66),.clk(clk),.wout(w101_66));
	PE pe101_67(.x(x67),.w(w101_66),.acc(r101_66),.res(r101_67),.clk(clk),.wout(w101_67));
	PE pe101_68(.x(x68),.w(w101_67),.acc(r101_67),.res(r101_68),.clk(clk),.wout(w101_68));
	PE pe101_69(.x(x69),.w(w101_68),.acc(r101_68),.res(r101_69),.clk(clk),.wout(w101_69));
	PE pe101_70(.x(x70),.w(w101_69),.acc(r101_69),.res(r101_70),.clk(clk),.wout(w101_70));
	PE pe101_71(.x(x71),.w(w101_70),.acc(r101_70),.res(r101_71),.clk(clk),.wout(w101_71));
	PE pe101_72(.x(x72),.w(w101_71),.acc(r101_71),.res(r101_72),.clk(clk),.wout(w101_72));
	PE pe101_73(.x(x73),.w(w101_72),.acc(r101_72),.res(r101_73),.clk(clk),.wout(w101_73));
	PE pe101_74(.x(x74),.w(w101_73),.acc(r101_73),.res(r101_74),.clk(clk),.wout(w101_74));
	PE pe101_75(.x(x75),.w(w101_74),.acc(r101_74),.res(r101_75),.clk(clk),.wout(w101_75));
	PE pe101_76(.x(x76),.w(w101_75),.acc(r101_75),.res(r101_76),.clk(clk),.wout(w101_76));
	PE pe101_77(.x(x77),.w(w101_76),.acc(r101_76),.res(r101_77),.clk(clk),.wout(w101_77));
	PE pe101_78(.x(x78),.w(w101_77),.acc(r101_77),.res(r101_78),.clk(clk),.wout(w101_78));
	PE pe101_79(.x(x79),.w(w101_78),.acc(r101_78),.res(r101_79),.clk(clk),.wout(w101_79));
	PE pe101_80(.x(x80),.w(w101_79),.acc(r101_79),.res(r101_80),.clk(clk),.wout(w101_80));
	PE pe101_81(.x(x81),.w(w101_80),.acc(r101_80),.res(r101_81),.clk(clk),.wout(w101_81));
	PE pe101_82(.x(x82),.w(w101_81),.acc(r101_81),.res(r101_82),.clk(clk),.wout(w101_82));
	PE pe101_83(.x(x83),.w(w101_82),.acc(r101_82),.res(r101_83),.clk(clk),.wout(w101_83));
	PE pe101_84(.x(x84),.w(w101_83),.acc(r101_83),.res(r101_84),.clk(clk),.wout(w101_84));
	PE pe101_85(.x(x85),.w(w101_84),.acc(r101_84),.res(r101_85),.clk(clk),.wout(w101_85));
	PE pe101_86(.x(x86),.w(w101_85),.acc(r101_85),.res(r101_86),.clk(clk),.wout(w101_86));
	PE pe101_87(.x(x87),.w(w101_86),.acc(r101_86),.res(r101_87),.clk(clk),.wout(w101_87));
	PE pe101_88(.x(x88),.w(w101_87),.acc(r101_87),.res(r101_88),.clk(clk),.wout(w101_88));
	PE pe101_89(.x(x89),.w(w101_88),.acc(r101_88),.res(r101_89),.clk(clk),.wout(w101_89));
	PE pe101_90(.x(x90),.w(w101_89),.acc(r101_89),.res(r101_90),.clk(clk),.wout(w101_90));
	PE pe101_91(.x(x91),.w(w101_90),.acc(r101_90),.res(r101_91),.clk(clk),.wout(w101_91));
	PE pe101_92(.x(x92),.w(w101_91),.acc(r101_91),.res(r101_92),.clk(clk),.wout(w101_92));
	PE pe101_93(.x(x93),.w(w101_92),.acc(r101_92),.res(r101_93),.clk(clk),.wout(w101_93));
	PE pe101_94(.x(x94),.w(w101_93),.acc(r101_93),.res(r101_94),.clk(clk),.wout(w101_94));
	PE pe101_95(.x(x95),.w(w101_94),.acc(r101_94),.res(r101_95),.clk(clk),.wout(w101_95));
	PE pe101_96(.x(x96),.w(w101_95),.acc(r101_95),.res(r101_96),.clk(clk),.wout(w101_96));
	PE pe101_97(.x(x97),.w(w101_96),.acc(r101_96),.res(r101_97),.clk(clk),.wout(w101_97));
	PE pe101_98(.x(x98),.w(w101_97),.acc(r101_97),.res(r101_98),.clk(clk),.wout(w101_98));
	PE pe101_99(.x(x99),.w(w101_98),.acc(r101_98),.res(r101_99),.clk(clk),.wout(w101_99));
	PE pe101_100(.x(x100),.w(w101_99),.acc(r101_99),.res(r101_100),.clk(clk),.wout(w101_100));
	PE pe101_101(.x(x101),.w(w101_100),.acc(r101_100),.res(r101_101),.clk(clk),.wout(w101_101));
	PE pe101_102(.x(x102),.w(w101_101),.acc(r101_101),.res(r101_102),.clk(clk),.wout(w101_102));
	PE pe101_103(.x(x103),.w(w101_102),.acc(r101_102),.res(r101_103),.clk(clk),.wout(w101_103));
	PE pe101_104(.x(x104),.w(w101_103),.acc(r101_103),.res(r101_104),.clk(clk),.wout(w101_104));
	PE pe101_105(.x(x105),.w(w101_104),.acc(r101_104),.res(r101_105),.clk(clk),.wout(w101_105));
	PE pe101_106(.x(x106),.w(w101_105),.acc(r101_105),.res(r101_106),.clk(clk),.wout(w101_106));
	PE pe101_107(.x(x107),.w(w101_106),.acc(r101_106),.res(r101_107),.clk(clk),.wout(w101_107));
	PE pe101_108(.x(x108),.w(w101_107),.acc(r101_107),.res(r101_108),.clk(clk),.wout(w101_108));
	PE pe101_109(.x(x109),.w(w101_108),.acc(r101_108),.res(r101_109),.clk(clk),.wout(w101_109));
	PE pe101_110(.x(x110),.w(w101_109),.acc(r101_109),.res(r101_110),.clk(clk),.wout(w101_110));
	PE pe101_111(.x(x111),.w(w101_110),.acc(r101_110),.res(r101_111),.clk(clk),.wout(w101_111));
	PE pe101_112(.x(x112),.w(w101_111),.acc(r101_111),.res(r101_112),.clk(clk),.wout(w101_112));
	PE pe101_113(.x(x113),.w(w101_112),.acc(r101_112),.res(r101_113),.clk(clk),.wout(w101_113));
	PE pe101_114(.x(x114),.w(w101_113),.acc(r101_113),.res(r101_114),.clk(clk),.wout(w101_114));
	PE pe101_115(.x(x115),.w(w101_114),.acc(r101_114),.res(r101_115),.clk(clk),.wout(w101_115));
	PE pe101_116(.x(x116),.w(w101_115),.acc(r101_115),.res(r101_116),.clk(clk),.wout(w101_116));
	PE pe101_117(.x(x117),.w(w101_116),.acc(r101_116),.res(r101_117),.clk(clk),.wout(w101_117));
	PE pe101_118(.x(x118),.w(w101_117),.acc(r101_117),.res(r101_118),.clk(clk),.wout(w101_118));
	PE pe101_119(.x(x119),.w(w101_118),.acc(r101_118),.res(r101_119),.clk(clk),.wout(w101_119));
	PE pe101_120(.x(x120),.w(w101_119),.acc(r101_119),.res(r101_120),.clk(clk),.wout(w101_120));
	PE pe101_121(.x(x121),.w(w101_120),.acc(r101_120),.res(r101_121),.clk(clk),.wout(w101_121));
	PE pe101_122(.x(x122),.w(w101_121),.acc(r101_121),.res(r101_122),.clk(clk),.wout(w101_122));
	PE pe101_123(.x(x123),.w(w101_122),.acc(r101_122),.res(r101_123),.clk(clk),.wout(w101_123));
	PE pe101_124(.x(x124),.w(w101_123),.acc(r101_123),.res(r101_124),.clk(clk),.wout(w101_124));
	PE pe101_125(.x(x125),.w(w101_124),.acc(r101_124),.res(r101_125),.clk(clk),.wout(w101_125));
	PE pe101_126(.x(x126),.w(w101_125),.acc(r101_125),.res(r101_126),.clk(clk),.wout(w101_126));
	PE pe101_127(.x(x127),.w(w101_126),.acc(r101_126),.res(result101),.clk(clk),.wout(weight101));

	PE pe102_0(.x(x0),.w(w102),.acc(32'h0),.res(r102_0),.clk(clk),.wout(w102_0));
	PE pe102_1(.x(x1),.w(w102_0),.acc(r102_0),.res(r102_1),.clk(clk),.wout(w102_1));
	PE pe102_2(.x(x2),.w(w102_1),.acc(r102_1),.res(r102_2),.clk(clk),.wout(w102_2));
	PE pe102_3(.x(x3),.w(w102_2),.acc(r102_2),.res(r102_3),.clk(clk),.wout(w102_3));
	PE pe102_4(.x(x4),.w(w102_3),.acc(r102_3),.res(r102_4),.clk(clk),.wout(w102_4));
	PE pe102_5(.x(x5),.w(w102_4),.acc(r102_4),.res(r102_5),.clk(clk),.wout(w102_5));
	PE pe102_6(.x(x6),.w(w102_5),.acc(r102_5),.res(r102_6),.clk(clk),.wout(w102_6));
	PE pe102_7(.x(x7),.w(w102_6),.acc(r102_6),.res(r102_7),.clk(clk),.wout(w102_7));
	PE pe102_8(.x(x8),.w(w102_7),.acc(r102_7),.res(r102_8),.clk(clk),.wout(w102_8));
	PE pe102_9(.x(x9),.w(w102_8),.acc(r102_8),.res(r102_9),.clk(clk),.wout(w102_9));
	PE pe102_10(.x(x10),.w(w102_9),.acc(r102_9),.res(r102_10),.clk(clk),.wout(w102_10));
	PE pe102_11(.x(x11),.w(w102_10),.acc(r102_10),.res(r102_11),.clk(clk),.wout(w102_11));
	PE pe102_12(.x(x12),.w(w102_11),.acc(r102_11),.res(r102_12),.clk(clk),.wout(w102_12));
	PE pe102_13(.x(x13),.w(w102_12),.acc(r102_12),.res(r102_13),.clk(clk),.wout(w102_13));
	PE pe102_14(.x(x14),.w(w102_13),.acc(r102_13),.res(r102_14),.clk(clk),.wout(w102_14));
	PE pe102_15(.x(x15),.w(w102_14),.acc(r102_14),.res(r102_15),.clk(clk),.wout(w102_15));
	PE pe102_16(.x(x16),.w(w102_15),.acc(r102_15),.res(r102_16),.clk(clk),.wout(w102_16));
	PE pe102_17(.x(x17),.w(w102_16),.acc(r102_16),.res(r102_17),.clk(clk),.wout(w102_17));
	PE pe102_18(.x(x18),.w(w102_17),.acc(r102_17),.res(r102_18),.clk(clk),.wout(w102_18));
	PE pe102_19(.x(x19),.w(w102_18),.acc(r102_18),.res(r102_19),.clk(clk),.wout(w102_19));
	PE pe102_20(.x(x20),.w(w102_19),.acc(r102_19),.res(r102_20),.clk(clk),.wout(w102_20));
	PE pe102_21(.x(x21),.w(w102_20),.acc(r102_20),.res(r102_21),.clk(clk),.wout(w102_21));
	PE pe102_22(.x(x22),.w(w102_21),.acc(r102_21),.res(r102_22),.clk(clk),.wout(w102_22));
	PE pe102_23(.x(x23),.w(w102_22),.acc(r102_22),.res(r102_23),.clk(clk),.wout(w102_23));
	PE pe102_24(.x(x24),.w(w102_23),.acc(r102_23),.res(r102_24),.clk(clk),.wout(w102_24));
	PE pe102_25(.x(x25),.w(w102_24),.acc(r102_24),.res(r102_25),.clk(clk),.wout(w102_25));
	PE pe102_26(.x(x26),.w(w102_25),.acc(r102_25),.res(r102_26),.clk(clk),.wout(w102_26));
	PE pe102_27(.x(x27),.w(w102_26),.acc(r102_26),.res(r102_27),.clk(clk),.wout(w102_27));
	PE pe102_28(.x(x28),.w(w102_27),.acc(r102_27),.res(r102_28),.clk(clk),.wout(w102_28));
	PE pe102_29(.x(x29),.w(w102_28),.acc(r102_28),.res(r102_29),.clk(clk),.wout(w102_29));
	PE pe102_30(.x(x30),.w(w102_29),.acc(r102_29),.res(r102_30),.clk(clk),.wout(w102_30));
	PE pe102_31(.x(x31),.w(w102_30),.acc(r102_30),.res(r102_31),.clk(clk),.wout(w102_31));
	PE pe102_32(.x(x32),.w(w102_31),.acc(r102_31),.res(r102_32),.clk(clk),.wout(w102_32));
	PE pe102_33(.x(x33),.w(w102_32),.acc(r102_32),.res(r102_33),.clk(clk),.wout(w102_33));
	PE pe102_34(.x(x34),.w(w102_33),.acc(r102_33),.res(r102_34),.clk(clk),.wout(w102_34));
	PE pe102_35(.x(x35),.w(w102_34),.acc(r102_34),.res(r102_35),.clk(clk),.wout(w102_35));
	PE pe102_36(.x(x36),.w(w102_35),.acc(r102_35),.res(r102_36),.clk(clk),.wout(w102_36));
	PE pe102_37(.x(x37),.w(w102_36),.acc(r102_36),.res(r102_37),.clk(clk),.wout(w102_37));
	PE pe102_38(.x(x38),.w(w102_37),.acc(r102_37),.res(r102_38),.clk(clk),.wout(w102_38));
	PE pe102_39(.x(x39),.w(w102_38),.acc(r102_38),.res(r102_39),.clk(clk),.wout(w102_39));
	PE pe102_40(.x(x40),.w(w102_39),.acc(r102_39),.res(r102_40),.clk(clk),.wout(w102_40));
	PE pe102_41(.x(x41),.w(w102_40),.acc(r102_40),.res(r102_41),.clk(clk),.wout(w102_41));
	PE pe102_42(.x(x42),.w(w102_41),.acc(r102_41),.res(r102_42),.clk(clk),.wout(w102_42));
	PE pe102_43(.x(x43),.w(w102_42),.acc(r102_42),.res(r102_43),.clk(clk),.wout(w102_43));
	PE pe102_44(.x(x44),.w(w102_43),.acc(r102_43),.res(r102_44),.clk(clk),.wout(w102_44));
	PE pe102_45(.x(x45),.w(w102_44),.acc(r102_44),.res(r102_45),.clk(clk),.wout(w102_45));
	PE pe102_46(.x(x46),.w(w102_45),.acc(r102_45),.res(r102_46),.clk(clk),.wout(w102_46));
	PE pe102_47(.x(x47),.w(w102_46),.acc(r102_46),.res(r102_47),.clk(clk),.wout(w102_47));
	PE pe102_48(.x(x48),.w(w102_47),.acc(r102_47),.res(r102_48),.clk(clk),.wout(w102_48));
	PE pe102_49(.x(x49),.w(w102_48),.acc(r102_48),.res(r102_49),.clk(clk),.wout(w102_49));
	PE pe102_50(.x(x50),.w(w102_49),.acc(r102_49),.res(r102_50),.clk(clk),.wout(w102_50));
	PE pe102_51(.x(x51),.w(w102_50),.acc(r102_50),.res(r102_51),.clk(clk),.wout(w102_51));
	PE pe102_52(.x(x52),.w(w102_51),.acc(r102_51),.res(r102_52),.clk(clk),.wout(w102_52));
	PE pe102_53(.x(x53),.w(w102_52),.acc(r102_52),.res(r102_53),.clk(clk),.wout(w102_53));
	PE pe102_54(.x(x54),.w(w102_53),.acc(r102_53),.res(r102_54),.clk(clk),.wout(w102_54));
	PE pe102_55(.x(x55),.w(w102_54),.acc(r102_54),.res(r102_55),.clk(clk),.wout(w102_55));
	PE pe102_56(.x(x56),.w(w102_55),.acc(r102_55),.res(r102_56),.clk(clk),.wout(w102_56));
	PE pe102_57(.x(x57),.w(w102_56),.acc(r102_56),.res(r102_57),.clk(clk),.wout(w102_57));
	PE pe102_58(.x(x58),.w(w102_57),.acc(r102_57),.res(r102_58),.clk(clk),.wout(w102_58));
	PE pe102_59(.x(x59),.w(w102_58),.acc(r102_58),.res(r102_59),.clk(clk),.wout(w102_59));
	PE pe102_60(.x(x60),.w(w102_59),.acc(r102_59),.res(r102_60),.clk(clk),.wout(w102_60));
	PE pe102_61(.x(x61),.w(w102_60),.acc(r102_60),.res(r102_61),.clk(clk),.wout(w102_61));
	PE pe102_62(.x(x62),.w(w102_61),.acc(r102_61),.res(r102_62),.clk(clk),.wout(w102_62));
	PE pe102_63(.x(x63),.w(w102_62),.acc(r102_62),.res(r102_63),.clk(clk),.wout(w102_63));
	PE pe102_64(.x(x64),.w(w102_63),.acc(r102_63),.res(r102_64),.clk(clk),.wout(w102_64));
	PE pe102_65(.x(x65),.w(w102_64),.acc(r102_64),.res(r102_65),.clk(clk),.wout(w102_65));
	PE pe102_66(.x(x66),.w(w102_65),.acc(r102_65),.res(r102_66),.clk(clk),.wout(w102_66));
	PE pe102_67(.x(x67),.w(w102_66),.acc(r102_66),.res(r102_67),.clk(clk),.wout(w102_67));
	PE pe102_68(.x(x68),.w(w102_67),.acc(r102_67),.res(r102_68),.clk(clk),.wout(w102_68));
	PE pe102_69(.x(x69),.w(w102_68),.acc(r102_68),.res(r102_69),.clk(clk),.wout(w102_69));
	PE pe102_70(.x(x70),.w(w102_69),.acc(r102_69),.res(r102_70),.clk(clk),.wout(w102_70));
	PE pe102_71(.x(x71),.w(w102_70),.acc(r102_70),.res(r102_71),.clk(clk),.wout(w102_71));
	PE pe102_72(.x(x72),.w(w102_71),.acc(r102_71),.res(r102_72),.clk(clk),.wout(w102_72));
	PE pe102_73(.x(x73),.w(w102_72),.acc(r102_72),.res(r102_73),.clk(clk),.wout(w102_73));
	PE pe102_74(.x(x74),.w(w102_73),.acc(r102_73),.res(r102_74),.clk(clk),.wout(w102_74));
	PE pe102_75(.x(x75),.w(w102_74),.acc(r102_74),.res(r102_75),.clk(clk),.wout(w102_75));
	PE pe102_76(.x(x76),.w(w102_75),.acc(r102_75),.res(r102_76),.clk(clk),.wout(w102_76));
	PE pe102_77(.x(x77),.w(w102_76),.acc(r102_76),.res(r102_77),.clk(clk),.wout(w102_77));
	PE pe102_78(.x(x78),.w(w102_77),.acc(r102_77),.res(r102_78),.clk(clk),.wout(w102_78));
	PE pe102_79(.x(x79),.w(w102_78),.acc(r102_78),.res(r102_79),.clk(clk),.wout(w102_79));
	PE pe102_80(.x(x80),.w(w102_79),.acc(r102_79),.res(r102_80),.clk(clk),.wout(w102_80));
	PE pe102_81(.x(x81),.w(w102_80),.acc(r102_80),.res(r102_81),.clk(clk),.wout(w102_81));
	PE pe102_82(.x(x82),.w(w102_81),.acc(r102_81),.res(r102_82),.clk(clk),.wout(w102_82));
	PE pe102_83(.x(x83),.w(w102_82),.acc(r102_82),.res(r102_83),.clk(clk),.wout(w102_83));
	PE pe102_84(.x(x84),.w(w102_83),.acc(r102_83),.res(r102_84),.clk(clk),.wout(w102_84));
	PE pe102_85(.x(x85),.w(w102_84),.acc(r102_84),.res(r102_85),.clk(clk),.wout(w102_85));
	PE pe102_86(.x(x86),.w(w102_85),.acc(r102_85),.res(r102_86),.clk(clk),.wout(w102_86));
	PE pe102_87(.x(x87),.w(w102_86),.acc(r102_86),.res(r102_87),.clk(clk),.wout(w102_87));
	PE pe102_88(.x(x88),.w(w102_87),.acc(r102_87),.res(r102_88),.clk(clk),.wout(w102_88));
	PE pe102_89(.x(x89),.w(w102_88),.acc(r102_88),.res(r102_89),.clk(clk),.wout(w102_89));
	PE pe102_90(.x(x90),.w(w102_89),.acc(r102_89),.res(r102_90),.clk(clk),.wout(w102_90));
	PE pe102_91(.x(x91),.w(w102_90),.acc(r102_90),.res(r102_91),.clk(clk),.wout(w102_91));
	PE pe102_92(.x(x92),.w(w102_91),.acc(r102_91),.res(r102_92),.clk(clk),.wout(w102_92));
	PE pe102_93(.x(x93),.w(w102_92),.acc(r102_92),.res(r102_93),.clk(clk),.wout(w102_93));
	PE pe102_94(.x(x94),.w(w102_93),.acc(r102_93),.res(r102_94),.clk(clk),.wout(w102_94));
	PE pe102_95(.x(x95),.w(w102_94),.acc(r102_94),.res(r102_95),.clk(clk),.wout(w102_95));
	PE pe102_96(.x(x96),.w(w102_95),.acc(r102_95),.res(r102_96),.clk(clk),.wout(w102_96));
	PE pe102_97(.x(x97),.w(w102_96),.acc(r102_96),.res(r102_97),.clk(clk),.wout(w102_97));
	PE pe102_98(.x(x98),.w(w102_97),.acc(r102_97),.res(r102_98),.clk(clk),.wout(w102_98));
	PE pe102_99(.x(x99),.w(w102_98),.acc(r102_98),.res(r102_99),.clk(clk),.wout(w102_99));
	PE pe102_100(.x(x100),.w(w102_99),.acc(r102_99),.res(r102_100),.clk(clk),.wout(w102_100));
	PE pe102_101(.x(x101),.w(w102_100),.acc(r102_100),.res(r102_101),.clk(clk),.wout(w102_101));
	PE pe102_102(.x(x102),.w(w102_101),.acc(r102_101),.res(r102_102),.clk(clk),.wout(w102_102));
	PE pe102_103(.x(x103),.w(w102_102),.acc(r102_102),.res(r102_103),.clk(clk),.wout(w102_103));
	PE pe102_104(.x(x104),.w(w102_103),.acc(r102_103),.res(r102_104),.clk(clk),.wout(w102_104));
	PE pe102_105(.x(x105),.w(w102_104),.acc(r102_104),.res(r102_105),.clk(clk),.wout(w102_105));
	PE pe102_106(.x(x106),.w(w102_105),.acc(r102_105),.res(r102_106),.clk(clk),.wout(w102_106));
	PE pe102_107(.x(x107),.w(w102_106),.acc(r102_106),.res(r102_107),.clk(clk),.wout(w102_107));
	PE pe102_108(.x(x108),.w(w102_107),.acc(r102_107),.res(r102_108),.clk(clk),.wout(w102_108));
	PE pe102_109(.x(x109),.w(w102_108),.acc(r102_108),.res(r102_109),.clk(clk),.wout(w102_109));
	PE pe102_110(.x(x110),.w(w102_109),.acc(r102_109),.res(r102_110),.clk(clk),.wout(w102_110));
	PE pe102_111(.x(x111),.w(w102_110),.acc(r102_110),.res(r102_111),.clk(clk),.wout(w102_111));
	PE pe102_112(.x(x112),.w(w102_111),.acc(r102_111),.res(r102_112),.clk(clk),.wout(w102_112));
	PE pe102_113(.x(x113),.w(w102_112),.acc(r102_112),.res(r102_113),.clk(clk),.wout(w102_113));
	PE pe102_114(.x(x114),.w(w102_113),.acc(r102_113),.res(r102_114),.clk(clk),.wout(w102_114));
	PE pe102_115(.x(x115),.w(w102_114),.acc(r102_114),.res(r102_115),.clk(clk),.wout(w102_115));
	PE pe102_116(.x(x116),.w(w102_115),.acc(r102_115),.res(r102_116),.clk(clk),.wout(w102_116));
	PE pe102_117(.x(x117),.w(w102_116),.acc(r102_116),.res(r102_117),.clk(clk),.wout(w102_117));
	PE pe102_118(.x(x118),.w(w102_117),.acc(r102_117),.res(r102_118),.clk(clk),.wout(w102_118));
	PE pe102_119(.x(x119),.w(w102_118),.acc(r102_118),.res(r102_119),.clk(clk),.wout(w102_119));
	PE pe102_120(.x(x120),.w(w102_119),.acc(r102_119),.res(r102_120),.clk(clk),.wout(w102_120));
	PE pe102_121(.x(x121),.w(w102_120),.acc(r102_120),.res(r102_121),.clk(clk),.wout(w102_121));
	PE pe102_122(.x(x122),.w(w102_121),.acc(r102_121),.res(r102_122),.clk(clk),.wout(w102_122));
	PE pe102_123(.x(x123),.w(w102_122),.acc(r102_122),.res(r102_123),.clk(clk),.wout(w102_123));
	PE pe102_124(.x(x124),.w(w102_123),.acc(r102_123),.res(r102_124),.clk(clk),.wout(w102_124));
	PE pe102_125(.x(x125),.w(w102_124),.acc(r102_124),.res(r102_125),.clk(clk),.wout(w102_125));
	PE pe102_126(.x(x126),.w(w102_125),.acc(r102_125),.res(r102_126),.clk(clk),.wout(w102_126));
	PE pe102_127(.x(x127),.w(w102_126),.acc(r102_126),.res(result102),.clk(clk),.wout(weight102));

	PE pe103_0(.x(x0),.w(w103),.acc(32'h0),.res(r103_0),.clk(clk),.wout(w103_0));
	PE pe103_1(.x(x1),.w(w103_0),.acc(r103_0),.res(r103_1),.clk(clk),.wout(w103_1));
	PE pe103_2(.x(x2),.w(w103_1),.acc(r103_1),.res(r103_2),.clk(clk),.wout(w103_2));
	PE pe103_3(.x(x3),.w(w103_2),.acc(r103_2),.res(r103_3),.clk(clk),.wout(w103_3));
	PE pe103_4(.x(x4),.w(w103_3),.acc(r103_3),.res(r103_4),.clk(clk),.wout(w103_4));
	PE pe103_5(.x(x5),.w(w103_4),.acc(r103_4),.res(r103_5),.clk(clk),.wout(w103_5));
	PE pe103_6(.x(x6),.w(w103_5),.acc(r103_5),.res(r103_6),.clk(clk),.wout(w103_6));
	PE pe103_7(.x(x7),.w(w103_6),.acc(r103_6),.res(r103_7),.clk(clk),.wout(w103_7));
	PE pe103_8(.x(x8),.w(w103_7),.acc(r103_7),.res(r103_8),.clk(clk),.wout(w103_8));
	PE pe103_9(.x(x9),.w(w103_8),.acc(r103_8),.res(r103_9),.clk(clk),.wout(w103_9));
	PE pe103_10(.x(x10),.w(w103_9),.acc(r103_9),.res(r103_10),.clk(clk),.wout(w103_10));
	PE pe103_11(.x(x11),.w(w103_10),.acc(r103_10),.res(r103_11),.clk(clk),.wout(w103_11));
	PE pe103_12(.x(x12),.w(w103_11),.acc(r103_11),.res(r103_12),.clk(clk),.wout(w103_12));
	PE pe103_13(.x(x13),.w(w103_12),.acc(r103_12),.res(r103_13),.clk(clk),.wout(w103_13));
	PE pe103_14(.x(x14),.w(w103_13),.acc(r103_13),.res(r103_14),.clk(clk),.wout(w103_14));
	PE pe103_15(.x(x15),.w(w103_14),.acc(r103_14),.res(r103_15),.clk(clk),.wout(w103_15));
	PE pe103_16(.x(x16),.w(w103_15),.acc(r103_15),.res(r103_16),.clk(clk),.wout(w103_16));
	PE pe103_17(.x(x17),.w(w103_16),.acc(r103_16),.res(r103_17),.clk(clk),.wout(w103_17));
	PE pe103_18(.x(x18),.w(w103_17),.acc(r103_17),.res(r103_18),.clk(clk),.wout(w103_18));
	PE pe103_19(.x(x19),.w(w103_18),.acc(r103_18),.res(r103_19),.clk(clk),.wout(w103_19));
	PE pe103_20(.x(x20),.w(w103_19),.acc(r103_19),.res(r103_20),.clk(clk),.wout(w103_20));
	PE pe103_21(.x(x21),.w(w103_20),.acc(r103_20),.res(r103_21),.clk(clk),.wout(w103_21));
	PE pe103_22(.x(x22),.w(w103_21),.acc(r103_21),.res(r103_22),.clk(clk),.wout(w103_22));
	PE pe103_23(.x(x23),.w(w103_22),.acc(r103_22),.res(r103_23),.clk(clk),.wout(w103_23));
	PE pe103_24(.x(x24),.w(w103_23),.acc(r103_23),.res(r103_24),.clk(clk),.wout(w103_24));
	PE pe103_25(.x(x25),.w(w103_24),.acc(r103_24),.res(r103_25),.clk(clk),.wout(w103_25));
	PE pe103_26(.x(x26),.w(w103_25),.acc(r103_25),.res(r103_26),.clk(clk),.wout(w103_26));
	PE pe103_27(.x(x27),.w(w103_26),.acc(r103_26),.res(r103_27),.clk(clk),.wout(w103_27));
	PE pe103_28(.x(x28),.w(w103_27),.acc(r103_27),.res(r103_28),.clk(clk),.wout(w103_28));
	PE pe103_29(.x(x29),.w(w103_28),.acc(r103_28),.res(r103_29),.clk(clk),.wout(w103_29));
	PE pe103_30(.x(x30),.w(w103_29),.acc(r103_29),.res(r103_30),.clk(clk),.wout(w103_30));
	PE pe103_31(.x(x31),.w(w103_30),.acc(r103_30),.res(r103_31),.clk(clk),.wout(w103_31));
	PE pe103_32(.x(x32),.w(w103_31),.acc(r103_31),.res(r103_32),.clk(clk),.wout(w103_32));
	PE pe103_33(.x(x33),.w(w103_32),.acc(r103_32),.res(r103_33),.clk(clk),.wout(w103_33));
	PE pe103_34(.x(x34),.w(w103_33),.acc(r103_33),.res(r103_34),.clk(clk),.wout(w103_34));
	PE pe103_35(.x(x35),.w(w103_34),.acc(r103_34),.res(r103_35),.clk(clk),.wout(w103_35));
	PE pe103_36(.x(x36),.w(w103_35),.acc(r103_35),.res(r103_36),.clk(clk),.wout(w103_36));
	PE pe103_37(.x(x37),.w(w103_36),.acc(r103_36),.res(r103_37),.clk(clk),.wout(w103_37));
	PE pe103_38(.x(x38),.w(w103_37),.acc(r103_37),.res(r103_38),.clk(clk),.wout(w103_38));
	PE pe103_39(.x(x39),.w(w103_38),.acc(r103_38),.res(r103_39),.clk(clk),.wout(w103_39));
	PE pe103_40(.x(x40),.w(w103_39),.acc(r103_39),.res(r103_40),.clk(clk),.wout(w103_40));
	PE pe103_41(.x(x41),.w(w103_40),.acc(r103_40),.res(r103_41),.clk(clk),.wout(w103_41));
	PE pe103_42(.x(x42),.w(w103_41),.acc(r103_41),.res(r103_42),.clk(clk),.wout(w103_42));
	PE pe103_43(.x(x43),.w(w103_42),.acc(r103_42),.res(r103_43),.clk(clk),.wout(w103_43));
	PE pe103_44(.x(x44),.w(w103_43),.acc(r103_43),.res(r103_44),.clk(clk),.wout(w103_44));
	PE pe103_45(.x(x45),.w(w103_44),.acc(r103_44),.res(r103_45),.clk(clk),.wout(w103_45));
	PE pe103_46(.x(x46),.w(w103_45),.acc(r103_45),.res(r103_46),.clk(clk),.wout(w103_46));
	PE pe103_47(.x(x47),.w(w103_46),.acc(r103_46),.res(r103_47),.clk(clk),.wout(w103_47));
	PE pe103_48(.x(x48),.w(w103_47),.acc(r103_47),.res(r103_48),.clk(clk),.wout(w103_48));
	PE pe103_49(.x(x49),.w(w103_48),.acc(r103_48),.res(r103_49),.clk(clk),.wout(w103_49));
	PE pe103_50(.x(x50),.w(w103_49),.acc(r103_49),.res(r103_50),.clk(clk),.wout(w103_50));
	PE pe103_51(.x(x51),.w(w103_50),.acc(r103_50),.res(r103_51),.clk(clk),.wout(w103_51));
	PE pe103_52(.x(x52),.w(w103_51),.acc(r103_51),.res(r103_52),.clk(clk),.wout(w103_52));
	PE pe103_53(.x(x53),.w(w103_52),.acc(r103_52),.res(r103_53),.clk(clk),.wout(w103_53));
	PE pe103_54(.x(x54),.w(w103_53),.acc(r103_53),.res(r103_54),.clk(clk),.wout(w103_54));
	PE pe103_55(.x(x55),.w(w103_54),.acc(r103_54),.res(r103_55),.clk(clk),.wout(w103_55));
	PE pe103_56(.x(x56),.w(w103_55),.acc(r103_55),.res(r103_56),.clk(clk),.wout(w103_56));
	PE pe103_57(.x(x57),.w(w103_56),.acc(r103_56),.res(r103_57),.clk(clk),.wout(w103_57));
	PE pe103_58(.x(x58),.w(w103_57),.acc(r103_57),.res(r103_58),.clk(clk),.wout(w103_58));
	PE pe103_59(.x(x59),.w(w103_58),.acc(r103_58),.res(r103_59),.clk(clk),.wout(w103_59));
	PE pe103_60(.x(x60),.w(w103_59),.acc(r103_59),.res(r103_60),.clk(clk),.wout(w103_60));
	PE pe103_61(.x(x61),.w(w103_60),.acc(r103_60),.res(r103_61),.clk(clk),.wout(w103_61));
	PE pe103_62(.x(x62),.w(w103_61),.acc(r103_61),.res(r103_62),.clk(clk),.wout(w103_62));
	PE pe103_63(.x(x63),.w(w103_62),.acc(r103_62),.res(r103_63),.clk(clk),.wout(w103_63));
	PE pe103_64(.x(x64),.w(w103_63),.acc(r103_63),.res(r103_64),.clk(clk),.wout(w103_64));
	PE pe103_65(.x(x65),.w(w103_64),.acc(r103_64),.res(r103_65),.clk(clk),.wout(w103_65));
	PE pe103_66(.x(x66),.w(w103_65),.acc(r103_65),.res(r103_66),.clk(clk),.wout(w103_66));
	PE pe103_67(.x(x67),.w(w103_66),.acc(r103_66),.res(r103_67),.clk(clk),.wout(w103_67));
	PE pe103_68(.x(x68),.w(w103_67),.acc(r103_67),.res(r103_68),.clk(clk),.wout(w103_68));
	PE pe103_69(.x(x69),.w(w103_68),.acc(r103_68),.res(r103_69),.clk(clk),.wout(w103_69));
	PE pe103_70(.x(x70),.w(w103_69),.acc(r103_69),.res(r103_70),.clk(clk),.wout(w103_70));
	PE pe103_71(.x(x71),.w(w103_70),.acc(r103_70),.res(r103_71),.clk(clk),.wout(w103_71));
	PE pe103_72(.x(x72),.w(w103_71),.acc(r103_71),.res(r103_72),.clk(clk),.wout(w103_72));
	PE pe103_73(.x(x73),.w(w103_72),.acc(r103_72),.res(r103_73),.clk(clk),.wout(w103_73));
	PE pe103_74(.x(x74),.w(w103_73),.acc(r103_73),.res(r103_74),.clk(clk),.wout(w103_74));
	PE pe103_75(.x(x75),.w(w103_74),.acc(r103_74),.res(r103_75),.clk(clk),.wout(w103_75));
	PE pe103_76(.x(x76),.w(w103_75),.acc(r103_75),.res(r103_76),.clk(clk),.wout(w103_76));
	PE pe103_77(.x(x77),.w(w103_76),.acc(r103_76),.res(r103_77),.clk(clk),.wout(w103_77));
	PE pe103_78(.x(x78),.w(w103_77),.acc(r103_77),.res(r103_78),.clk(clk),.wout(w103_78));
	PE pe103_79(.x(x79),.w(w103_78),.acc(r103_78),.res(r103_79),.clk(clk),.wout(w103_79));
	PE pe103_80(.x(x80),.w(w103_79),.acc(r103_79),.res(r103_80),.clk(clk),.wout(w103_80));
	PE pe103_81(.x(x81),.w(w103_80),.acc(r103_80),.res(r103_81),.clk(clk),.wout(w103_81));
	PE pe103_82(.x(x82),.w(w103_81),.acc(r103_81),.res(r103_82),.clk(clk),.wout(w103_82));
	PE pe103_83(.x(x83),.w(w103_82),.acc(r103_82),.res(r103_83),.clk(clk),.wout(w103_83));
	PE pe103_84(.x(x84),.w(w103_83),.acc(r103_83),.res(r103_84),.clk(clk),.wout(w103_84));
	PE pe103_85(.x(x85),.w(w103_84),.acc(r103_84),.res(r103_85),.clk(clk),.wout(w103_85));
	PE pe103_86(.x(x86),.w(w103_85),.acc(r103_85),.res(r103_86),.clk(clk),.wout(w103_86));
	PE pe103_87(.x(x87),.w(w103_86),.acc(r103_86),.res(r103_87),.clk(clk),.wout(w103_87));
	PE pe103_88(.x(x88),.w(w103_87),.acc(r103_87),.res(r103_88),.clk(clk),.wout(w103_88));
	PE pe103_89(.x(x89),.w(w103_88),.acc(r103_88),.res(r103_89),.clk(clk),.wout(w103_89));
	PE pe103_90(.x(x90),.w(w103_89),.acc(r103_89),.res(r103_90),.clk(clk),.wout(w103_90));
	PE pe103_91(.x(x91),.w(w103_90),.acc(r103_90),.res(r103_91),.clk(clk),.wout(w103_91));
	PE pe103_92(.x(x92),.w(w103_91),.acc(r103_91),.res(r103_92),.clk(clk),.wout(w103_92));
	PE pe103_93(.x(x93),.w(w103_92),.acc(r103_92),.res(r103_93),.clk(clk),.wout(w103_93));
	PE pe103_94(.x(x94),.w(w103_93),.acc(r103_93),.res(r103_94),.clk(clk),.wout(w103_94));
	PE pe103_95(.x(x95),.w(w103_94),.acc(r103_94),.res(r103_95),.clk(clk),.wout(w103_95));
	PE pe103_96(.x(x96),.w(w103_95),.acc(r103_95),.res(r103_96),.clk(clk),.wout(w103_96));
	PE pe103_97(.x(x97),.w(w103_96),.acc(r103_96),.res(r103_97),.clk(clk),.wout(w103_97));
	PE pe103_98(.x(x98),.w(w103_97),.acc(r103_97),.res(r103_98),.clk(clk),.wout(w103_98));
	PE pe103_99(.x(x99),.w(w103_98),.acc(r103_98),.res(r103_99),.clk(clk),.wout(w103_99));
	PE pe103_100(.x(x100),.w(w103_99),.acc(r103_99),.res(r103_100),.clk(clk),.wout(w103_100));
	PE pe103_101(.x(x101),.w(w103_100),.acc(r103_100),.res(r103_101),.clk(clk),.wout(w103_101));
	PE pe103_102(.x(x102),.w(w103_101),.acc(r103_101),.res(r103_102),.clk(clk),.wout(w103_102));
	PE pe103_103(.x(x103),.w(w103_102),.acc(r103_102),.res(r103_103),.clk(clk),.wout(w103_103));
	PE pe103_104(.x(x104),.w(w103_103),.acc(r103_103),.res(r103_104),.clk(clk),.wout(w103_104));
	PE pe103_105(.x(x105),.w(w103_104),.acc(r103_104),.res(r103_105),.clk(clk),.wout(w103_105));
	PE pe103_106(.x(x106),.w(w103_105),.acc(r103_105),.res(r103_106),.clk(clk),.wout(w103_106));
	PE pe103_107(.x(x107),.w(w103_106),.acc(r103_106),.res(r103_107),.clk(clk),.wout(w103_107));
	PE pe103_108(.x(x108),.w(w103_107),.acc(r103_107),.res(r103_108),.clk(clk),.wout(w103_108));
	PE pe103_109(.x(x109),.w(w103_108),.acc(r103_108),.res(r103_109),.clk(clk),.wout(w103_109));
	PE pe103_110(.x(x110),.w(w103_109),.acc(r103_109),.res(r103_110),.clk(clk),.wout(w103_110));
	PE pe103_111(.x(x111),.w(w103_110),.acc(r103_110),.res(r103_111),.clk(clk),.wout(w103_111));
	PE pe103_112(.x(x112),.w(w103_111),.acc(r103_111),.res(r103_112),.clk(clk),.wout(w103_112));
	PE pe103_113(.x(x113),.w(w103_112),.acc(r103_112),.res(r103_113),.clk(clk),.wout(w103_113));
	PE pe103_114(.x(x114),.w(w103_113),.acc(r103_113),.res(r103_114),.clk(clk),.wout(w103_114));
	PE pe103_115(.x(x115),.w(w103_114),.acc(r103_114),.res(r103_115),.clk(clk),.wout(w103_115));
	PE pe103_116(.x(x116),.w(w103_115),.acc(r103_115),.res(r103_116),.clk(clk),.wout(w103_116));
	PE pe103_117(.x(x117),.w(w103_116),.acc(r103_116),.res(r103_117),.clk(clk),.wout(w103_117));
	PE pe103_118(.x(x118),.w(w103_117),.acc(r103_117),.res(r103_118),.clk(clk),.wout(w103_118));
	PE pe103_119(.x(x119),.w(w103_118),.acc(r103_118),.res(r103_119),.clk(clk),.wout(w103_119));
	PE pe103_120(.x(x120),.w(w103_119),.acc(r103_119),.res(r103_120),.clk(clk),.wout(w103_120));
	PE pe103_121(.x(x121),.w(w103_120),.acc(r103_120),.res(r103_121),.clk(clk),.wout(w103_121));
	PE pe103_122(.x(x122),.w(w103_121),.acc(r103_121),.res(r103_122),.clk(clk),.wout(w103_122));
	PE pe103_123(.x(x123),.w(w103_122),.acc(r103_122),.res(r103_123),.clk(clk),.wout(w103_123));
	PE pe103_124(.x(x124),.w(w103_123),.acc(r103_123),.res(r103_124),.clk(clk),.wout(w103_124));
	PE pe103_125(.x(x125),.w(w103_124),.acc(r103_124),.res(r103_125),.clk(clk),.wout(w103_125));
	PE pe103_126(.x(x126),.w(w103_125),.acc(r103_125),.res(r103_126),.clk(clk),.wout(w103_126));
	PE pe103_127(.x(x127),.w(w103_126),.acc(r103_126),.res(result103),.clk(clk),.wout(weight103));

	PE pe104_0(.x(x0),.w(w104),.acc(32'h0),.res(r104_0),.clk(clk),.wout(w104_0));
	PE pe104_1(.x(x1),.w(w104_0),.acc(r104_0),.res(r104_1),.clk(clk),.wout(w104_1));
	PE pe104_2(.x(x2),.w(w104_1),.acc(r104_1),.res(r104_2),.clk(clk),.wout(w104_2));
	PE pe104_3(.x(x3),.w(w104_2),.acc(r104_2),.res(r104_3),.clk(clk),.wout(w104_3));
	PE pe104_4(.x(x4),.w(w104_3),.acc(r104_3),.res(r104_4),.clk(clk),.wout(w104_4));
	PE pe104_5(.x(x5),.w(w104_4),.acc(r104_4),.res(r104_5),.clk(clk),.wout(w104_5));
	PE pe104_6(.x(x6),.w(w104_5),.acc(r104_5),.res(r104_6),.clk(clk),.wout(w104_6));
	PE pe104_7(.x(x7),.w(w104_6),.acc(r104_6),.res(r104_7),.clk(clk),.wout(w104_7));
	PE pe104_8(.x(x8),.w(w104_7),.acc(r104_7),.res(r104_8),.clk(clk),.wout(w104_8));
	PE pe104_9(.x(x9),.w(w104_8),.acc(r104_8),.res(r104_9),.clk(clk),.wout(w104_9));
	PE pe104_10(.x(x10),.w(w104_9),.acc(r104_9),.res(r104_10),.clk(clk),.wout(w104_10));
	PE pe104_11(.x(x11),.w(w104_10),.acc(r104_10),.res(r104_11),.clk(clk),.wout(w104_11));
	PE pe104_12(.x(x12),.w(w104_11),.acc(r104_11),.res(r104_12),.clk(clk),.wout(w104_12));
	PE pe104_13(.x(x13),.w(w104_12),.acc(r104_12),.res(r104_13),.clk(clk),.wout(w104_13));
	PE pe104_14(.x(x14),.w(w104_13),.acc(r104_13),.res(r104_14),.clk(clk),.wout(w104_14));
	PE pe104_15(.x(x15),.w(w104_14),.acc(r104_14),.res(r104_15),.clk(clk),.wout(w104_15));
	PE pe104_16(.x(x16),.w(w104_15),.acc(r104_15),.res(r104_16),.clk(clk),.wout(w104_16));
	PE pe104_17(.x(x17),.w(w104_16),.acc(r104_16),.res(r104_17),.clk(clk),.wout(w104_17));
	PE pe104_18(.x(x18),.w(w104_17),.acc(r104_17),.res(r104_18),.clk(clk),.wout(w104_18));
	PE pe104_19(.x(x19),.w(w104_18),.acc(r104_18),.res(r104_19),.clk(clk),.wout(w104_19));
	PE pe104_20(.x(x20),.w(w104_19),.acc(r104_19),.res(r104_20),.clk(clk),.wout(w104_20));
	PE pe104_21(.x(x21),.w(w104_20),.acc(r104_20),.res(r104_21),.clk(clk),.wout(w104_21));
	PE pe104_22(.x(x22),.w(w104_21),.acc(r104_21),.res(r104_22),.clk(clk),.wout(w104_22));
	PE pe104_23(.x(x23),.w(w104_22),.acc(r104_22),.res(r104_23),.clk(clk),.wout(w104_23));
	PE pe104_24(.x(x24),.w(w104_23),.acc(r104_23),.res(r104_24),.clk(clk),.wout(w104_24));
	PE pe104_25(.x(x25),.w(w104_24),.acc(r104_24),.res(r104_25),.clk(clk),.wout(w104_25));
	PE pe104_26(.x(x26),.w(w104_25),.acc(r104_25),.res(r104_26),.clk(clk),.wout(w104_26));
	PE pe104_27(.x(x27),.w(w104_26),.acc(r104_26),.res(r104_27),.clk(clk),.wout(w104_27));
	PE pe104_28(.x(x28),.w(w104_27),.acc(r104_27),.res(r104_28),.clk(clk),.wout(w104_28));
	PE pe104_29(.x(x29),.w(w104_28),.acc(r104_28),.res(r104_29),.clk(clk),.wout(w104_29));
	PE pe104_30(.x(x30),.w(w104_29),.acc(r104_29),.res(r104_30),.clk(clk),.wout(w104_30));
	PE pe104_31(.x(x31),.w(w104_30),.acc(r104_30),.res(r104_31),.clk(clk),.wout(w104_31));
	PE pe104_32(.x(x32),.w(w104_31),.acc(r104_31),.res(r104_32),.clk(clk),.wout(w104_32));
	PE pe104_33(.x(x33),.w(w104_32),.acc(r104_32),.res(r104_33),.clk(clk),.wout(w104_33));
	PE pe104_34(.x(x34),.w(w104_33),.acc(r104_33),.res(r104_34),.clk(clk),.wout(w104_34));
	PE pe104_35(.x(x35),.w(w104_34),.acc(r104_34),.res(r104_35),.clk(clk),.wout(w104_35));
	PE pe104_36(.x(x36),.w(w104_35),.acc(r104_35),.res(r104_36),.clk(clk),.wout(w104_36));
	PE pe104_37(.x(x37),.w(w104_36),.acc(r104_36),.res(r104_37),.clk(clk),.wout(w104_37));
	PE pe104_38(.x(x38),.w(w104_37),.acc(r104_37),.res(r104_38),.clk(clk),.wout(w104_38));
	PE pe104_39(.x(x39),.w(w104_38),.acc(r104_38),.res(r104_39),.clk(clk),.wout(w104_39));
	PE pe104_40(.x(x40),.w(w104_39),.acc(r104_39),.res(r104_40),.clk(clk),.wout(w104_40));
	PE pe104_41(.x(x41),.w(w104_40),.acc(r104_40),.res(r104_41),.clk(clk),.wout(w104_41));
	PE pe104_42(.x(x42),.w(w104_41),.acc(r104_41),.res(r104_42),.clk(clk),.wout(w104_42));
	PE pe104_43(.x(x43),.w(w104_42),.acc(r104_42),.res(r104_43),.clk(clk),.wout(w104_43));
	PE pe104_44(.x(x44),.w(w104_43),.acc(r104_43),.res(r104_44),.clk(clk),.wout(w104_44));
	PE pe104_45(.x(x45),.w(w104_44),.acc(r104_44),.res(r104_45),.clk(clk),.wout(w104_45));
	PE pe104_46(.x(x46),.w(w104_45),.acc(r104_45),.res(r104_46),.clk(clk),.wout(w104_46));
	PE pe104_47(.x(x47),.w(w104_46),.acc(r104_46),.res(r104_47),.clk(clk),.wout(w104_47));
	PE pe104_48(.x(x48),.w(w104_47),.acc(r104_47),.res(r104_48),.clk(clk),.wout(w104_48));
	PE pe104_49(.x(x49),.w(w104_48),.acc(r104_48),.res(r104_49),.clk(clk),.wout(w104_49));
	PE pe104_50(.x(x50),.w(w104_49),.acc(r104_49),.res(r104_50),.clk(clk),.wout(w104_50));
	PE pe104_51(.x(x51),.w(w104_50),.acc(r104_50),.res(r104_51),.clk(clk),.wout(w104_51));
	PE pe104_52(.x(x52),.w(w104_51),.acc(r104_51),.res(r104_52),.clk(clk),.wout(w104_52));
	PE pe104_53(.x(x53),.w(w104_52),.acc(r104_52),.res(r104_53),.clk(clk),.wout(w104_53));
	PE pe104_54(.x(x54),.w(w104_53),.acc(r104_53),.res(r104_54),.clk(clk),.wout(w104_54));
	PE pe104_55(.x(x55),.w(w104_54),.acc(r104_54),.res(r104_55),.clk(clk),.wout(w104_55));
	PE pe104_56(.x(x56),.w(w104_55),.acc(r104_55),.res(r104_56),.clk(clk),.wout(w104_56));
	PE pe104_57(.x(x57),.w(w104_56),.acc(r104_56),.res(r104_57),.clk(clk),.wout(w104_57));
	PE pe104_58(.x(x58),.w(w104_57),.acc(r104_57),.res(r104_58),.clk(clk),.wout(w104_58));
	PE pe104_59(.x(x59),.w(w104_58),.acc(r104_58),.res(r104_59),.clk(clk),.wout(w104_59));
	PE pe104_60(.x(x60),.w(w104_59),.acc(r104_59),.res(r104_60),.clk(clk),.wout(w104_60));
	PE pe104_61(.x(x61),.w(w104_60),.acc(r104_60),.res(r104_61),.clk(clk),.wout(w104_61));
	PE pe104_62(.x(x62),.w(w104_61),.acc(r104_61),.res(r104_62),.clk(clk),.wout(w104_62));
	PE pe104_63(.x(x63),.w(w104_62),.acc(r104_62),.res(r104_63),.clk(clk),.wout(w104_63));
	PE pe104_64(.x(x64),.w(w104_63),.acc(r104_63),.res(r104_64),.clk(clk),.wout(w104_64));
	PE pe104_65(.x(x65),.w(w104_64),.acc(r104_64),.res(r104_65),.clk(clk),.wout(w104_65));
	PE pe104_66(.x(x66),.w(w104_65),.acc(r104_65),.res(r104_66),.clk(clk),.wout(w104_66));
	PE pe104_67(.x(x67),.w(w104_66),.acc(r104_66),.res(r104_67),.clk(clk),.wout(w104_67));
	PE pe104_68(.x(x68),.w(w104_67),.acc(r104_67),.res(r104_68),.clk(clk),.wout(w104_68));
	PE pe104_69(.x(x69),.w(w104_68),.acc(r104_68),.res(r104_69),.clk(clk),.wout(w104_69));
	PE pe104_70(.x(x70),.w(w104_69),.acc(r104_69),.res(r104_70),.clk(clk),.wout(w104_70));
	PE pe104_71(.x(x71),.w(w104_70),.acc(r104_70),.res(r104_71),.clk(clk),.wout(w104_71));
	PE pe104_72(.x(x72),.w(w104_71),.acc(r104_71),.res(r104_72),.clk(clk),.wout(w104_72));
	PE pe104_73(.x(x73),.w(w104_72),.acc(r104_72),.res(r104_73),.clk(clk),.wout(w104_73));
	PE pe104_74(.x(x74),.w(w104_73),.acc(r104_73),.res(r104_74),.clk(clk),.wout(w104_74));
	PE pe104_75(.x(x75),.w(w104_74),.acc(r104_74),.res(r104_75),.clk(clk),.wout(w104_75));
	PE pe104_76(.x(x76),.w(w104_75),.acc(r104_75),.res(r104_76),.clk(clk),.wout(w104_76));
	PE pe104_77(.x(x77),.w(w104_76),.acc(r104_76),.res(r104_77),.clk(clk),.wout(w104_77));
	PE pe104_78(.x(x78),.w(w104_77),.acc(r104_77),.res(r104_78),.clk(clk),.wout(w104_78));
	PE pe104_79(.x(x79),.w(w104_78),.acc(r104_78),.res(r104_79),.clk(clk),.wout(w104_79));
	PE pe104_80(.x(x80),.w(w104_79),.acc(r104_79),.res(r104_80),.clk(clk),.wout(w104_80));
	PE pe104_81(.x(x81),.w(w104_80),.acc(r104_80),.res(r104_81),.clk(clk),.wout(w104_81));
	PE pe104_82(.x(x82),.w(w104_81),.acc(r104_81),.res(r104_82),.clk(clk),.wout(w104_82));
	PE pe104_83(.x(x83),.w(w104_82),.acc(r104_82),.res(r104_83),.clk(clk),.wout(w104_83));
	PE pe104_84(.x(x84),.w(w104_83),.acc(r104_83),.res(r104_84),.clk(clk),.wout(w104_84));
	PE pe104_85(.x(x85),.w(w104_84),.acc(r104_84),.res(r104_85),.clk(clk),.wout(w104_85));
	PE pe104_86(.x(x86),.w(w104_85),.acc(r104_85),.res(r104_86),.clk(clk),.wout(w104_86));
	PE pe104_87(.x(x87),.w(w104_86),.acc(r104_86),.res(r104_87),.clk(clk),.wout(w104_87));
	PE pe104_88(.x(x88),.w(w104_87),.acc(r104_87),.res(r104_88),.clk(clk),.wout(w104_88));
	PE pe104_89(.x(x89),.w(w104_88),.acc(r104_88),.res(r104_89),.clk(clk),.wout(w104_89));
	PE pe104_90(.x(x90),.w(w104_89),.acc(r104_89),.res(r104_90),.clk(clk),.wout(w104_90));
	PE pe104_91(.x(x91),.w(w104_90),.acc(r104_90),.res(r104_91),.clk(clk),.wout(w104_91));
	PE pe104_92(.x(x92),.w(w104_91),.acc(r104_91),.res(r104_92),.clk(clk),.wout(w104_92));
	PE pe104_93(.x(x93),.w(w104_92),.acc(r104_92),.res(r104_93),.clk(clk),.wout(w104_93));
	PE pe104_94(.x(x94),.w(w104_93),.acc(r104_93),.res(r104_94),.clk(clk),.wout(w104_94));
	PE pe104_95(.x(x95),.w(w104_94),.acc(r104_94),.res(r104_95),.clk(clk),.wout(w104_95));
	PE pe104_96(.x(x96),.w(w104_95),.acc(r104_95),.res(r104_96),.clk(clk),.wout(w104_96));
	PE pe104_97(.x(x97),.w(w104_96),.acc(r104_96),.res(r104_97),.clk(clk),.wout(w104_97));
	PE pe104_98(.x(x98),.w(w104_97),.acc(r104_97),.res(r104_98),.clk(clk),.wout(w104_98));
	PE pe104_99(.x(x99),.w(w104_98),.acc(r104_98),.res(r104_99),.clk(clk),.wout(w104_99));
	PE pe104_100(.x(x100),.w(w104_99),.acc(r104_99),.res(r104_100),.clk(clk),.wout(w104_100));
	PE pe104_101(.x(x101),.w(w104_100),.acc(r104_100),.res(r104_101),.clk(clk),.wout(w104_101));
	PE pe104_102(.x(x102),.w(w104_101),.acc(r104_101),.res(r104_102),.clk(clk),.wout(w104_102));
	PE pe104_103(.x(x103),.w(w104_102),.acc(r104_102),.res(r104_103),.clk(clk),.wout(w104_103));
	PE pe104_104(.x(x104),.w(w104_103),.acc(r104_103),.res(r104_104),.clk(clk),.wout(w104_104));
	PE pe104_105(.x(x105),.w(w104_104),.acc(r104_104),.res(r104_105),.clk(clk),.wout(w104_105));
	PE pe104_106(.x(x106),.w(w104_105),.acc(r104_105),.res(r104_106),.clk(clk),.wout(w104_106));
	PE pe104_107(.x(x107),.w(w104_106),.acc(r104_106),.res(r104_107),.clk(clk),.wout(w104_107));
	PE pe104_108(.x(x108),.w(w104_107),.acc(r104_107),.res(r104_108),.clk(clk),.wout(w104_108));
	PE pe104_109(.x(x109),.w(w104_108),.acc(r104_108),.res(r104_109),.clk(clk),.wout(w104_109));
	PE pe104_110(.x(x110),.w(w104_109),.acc(r104_109),.res(r104_110),.clk(clk),.wout(w104_110));
	PE pe104_111(.x(x111),.w(w104_110),.acc(r104_110),.res(r104_111),.clk(clk),.wout(w104_111));
	PE pe104_112(.x(x112),.w(w104_111),.acc(r104_111),.res(r104_112),.clk(clk),.wout(w104_112));
	PE pe104_113(.x(x113),.w(w104_112),.acc(r104_112),.res(r104_113),.clk(clk),.wout(w104_113));
	PE pe104_114(.x(x114),.w(w104_113),.acc(r104_113),.res(r104_114),.clk(clk),.wout(w104_114));
	PE pe104_115(.x(x115),.w(w104_114),.acc(r104_114),.res(r104_115),.clk(clk),.wout(w104_115));
	PE pe104_116(.x(x116),.w(w104_115),.acc(r104_115),.res(r104_116),.clk(clk),.wout(w104_116));
	PE pe104_117(.x(x117),.w(w104_116),.acc(r104_116),.res(r104_117),.clk(clk),.wout(w104_117));
	PE pe104_118(.x(x118),.w(w104_117),.acc(r104_117),.res(r104_118),.clk(clk),.wout(w104_118));
	PE pe104_119(.x(x119),.w(w104_118),.acc(r104_118),.res(r104_119),.clk(clk),.wout(w104_119));
	PE pe104_120(.x(x120),.w(w104_119),.acc(r104_119),.res(r104_120),.clk(clk),.wout(w104_120));
	PE pe104_121(.x(x121),.w(w104_120),.acc(r104_120),.res(r104_121),.clk(clk),.wout(w104_121));
	PE pe104_122(.x(x122),.w(w104_121),.acc(r104_121),.res(r104_122),.clk(clk),.wout(w104_122));
	PE pe104_123(.x(x123),.w(w104_122),.acc(r104_122),.res(r104_123),.clk(clk),.wout(w104_123));
	PE pe104_124(.x(x124),.w(w104_123),.acc(r104_123),.res(r104_124),.clk(clk),.wout(w104_124));
	PE pe104_125(.x(x125),.w(w104_124),.acc(r104_124),.res(r104_125),.clk(clk),.wout(w104_125));
	PE pe104_126(.x(x126),.w(w104_125),.acc(r104_125),.res(r104_126),.clk(clk),.wout(w104_126));
	PE pe104_127(.x(x127),.w(w104_126),.acc(r104_126),.res(result104),.clk(clk),.wout(weight104));

	PE pe105_0(.x(x0),.w(w105),.acc(32'h0),.res(r105_0),.clk(clk),.wout(w105_0));
	PE pe105_1(.x(x1),.w(w105_0),.acc(r105_0),.res(r105_1),.clk(clk),.wout(w105_1));
	PE pe105_2(.x(x2),.w(w105_1),.acc(r105_1),.res(r105_2),.clk(clk),.wout(w105_2));
	PE pe105_3(.x(x3),.w(w105_2),.acc(r105_2),.res(r105_3),.clk(clk),.wout(w105_3));
	PE pe105_4(.x(x4),.w(w105_3),.acc(r105_3),.res(r105_4),.clk(clk),.wout(w105_4));
	PE pe105_5(.x(x5),.w(w105_4),.acc(r105_4),.res(r105_5),.clk(clk),.wout(w105_5));
	PE pe105_6(.x(x6),.w(w105_5),.acc(r105_5),.res(r105_6),.clk(clk),.wout(w105_6));
	PE pe105_7(.x(x7),.w(w105_6),.acc(r105_6),.res(r105_7),.clk(clk),.wout(w105_7));
	PE pe105_8(.x(x8),.w(w105_7),.acc(r105_7),.res(r105_8),.clk(clk),.wout(w105_8));
	PE pe105_9(.x(x9),.w(w105_8),.acc(r105_8),.res(r105_9),.clk(clk),.wout(w105_9));
	PE pe105_10(.x(x10),.w(w105_9),.acc(r105_9),.res(r105_10),.clk(clk),.wout(w105_10));
	PE pe105_11(.x(x11),.w(w105_10),.acc(r105_10),.res(r105_11),.clk(clk),.wout(w105_11));
	PE pe105_12(.x(x12),.w(w105_11),.acc(r105_11),.res(r105_12),.clk(clk),.wout(w105_12));
	PE pe105_13(.x(x13),.w(w105_12),.acc(r105_12),.res(r105_13),.clk(clk),.wout(w105_13));
	PE pe105_14(.x(x14),.w(w105_13),.acc(r105_13),.res(r105_14),.clk(clk),.wout(w105_14));
	PE pe105_15(.x(x15),.w(w105_14),.acc(r105_14),.res(r105_15),.clk(clk),.wout(w105_15));
	PE pe105_16(.x(x16),.w(w105_15),.acc(r105_15),.res(r105_16),.clk(clk),.wout(w105_16));
	PE pe105_17(.x(x17),.w(w105_16),.acc(r105_16),.res(r105_17),.clk(clk),.wout(w105_17));
	PE pe105_18(.x(x18),.w(w105_17),.acc(r105_17),.res(r105_18),.clk(clk),.wout(w105_18));
	PE pe105_19(.x(x19),.w(w105_18),.acc(r105_18),.res(r105_19),.clk(clk),.wout(w105_19));
	PE pe105_20(.x(x20),.w(w105_19),.acc(r105_19),.res(r105_20),.clk(clk),.wout(w105_20));
	PE pe105_21(.x(x21),.w(w105_20),.acc(r105_20),.res(r105_21),.clk(clk),.wout(w105_21));
	PE pe105_22(.x(x22),.w(w105_21),.acc(r105_21),.res(r105_22),.clk(clk),.wout(w105_22));
	PE pe105_23(.x(x23),.w(w105_22),.acc(r105_22),.res(r105_23),.clk(clk),.wout(w105_23));
	PE pe105_24(.x(x24),.w(w105_23),.acc(r105_23),.res(r105_24),.clk(clk),.wout(w105_24));
	PE pe105_25(.x(x25),.w(w105_24),.acc(r105_24),.res(r105_25),.clk(clk),.wout(w105_25));
	PE pe105_26(.x(x26),.w(w105_25),.acc(r105_25),.res(r105_26),.clk(clk),.wout(w105_26));
	PE pe105_27(.x(x27),.w(w105_26),.acc(r105_26),.res(r105_27),.clk(clk),.wout(w105_27));
	PE pe105_28(.x(x28),.w(w105_27),.acc(r105_27),.res(r105_28),.clk(clk),.wout(w105_28));
	PE pe105_29(.x(x29),.w(w105_28),.acc(r105_28),.res(r105_29),.clk(clk),.wout(w105_29));
	PE pe105_30(.x(x30),.w(w105_29),.acc(r105_29),.res(r105_30),.clk(clk),.wout(w105_30));
	PE pe105_31(.x(x31),.w(w105_30),.acc(r105_30),.res(r105_31),.clk(clk),.wout(w105_31));
	PE pe105_32(.x(x32),.w(w105_31),.acc(r105_31),.res(r105_32),.clk(clk),.wout(w105_32));
	PE pe105_33(.x(x33),.w(w105_32),.acc(r105_32),.res(r105_33),.clk(clk),.wout(w105_33));
	PE pe105_34(.x(x34),.w(w105_33),.acc(r105_33),.res(r105_34),.clk(clk),.wout(w105_34));
	PE pe105_35(.x(x35),.w(w105_34),.acc(r105_34),.res(r105_35),.clk(clk),.wout(w105_35));
	PE pe105_36(.x(x36),.w(w105_35),.acc(r105_35),.res(r105_36),.clk(clk),.wout(w105_36));
	PE pe105_37(.x(x37),.w(w105_36),.acc(r105_36),.res(r105_37),.clk(clk),.wout(w105_37));
	PE pe105_38(.x(x38),.w(w105_37),.acc(r105_37),.res(r105_38),.clk(clk),.wout(w105_38));
	PE pe105_39(.x(x39),.w(w105_38),.acc(r105_38),.res(r105_39),.clk(clk),.wout(w105_39));
	PE pe105_40(.x(x40),.w(w105_39),.acc(r105_39),.res(r105_40),.clk(clk),.wout(w105_40));
	PE pe105_41(.x(x41),.w(w105_40),.acc(r105_40),.res(r105_41),.clk(clk),.wout(w105_41));
	PE pe105_42(.x(x42),.w(w105_41),.acc(r105_41),.res(r105_42),.clk(clk),.wout(w105_42));
	PE pe105_43(.x(x43),.w(w105_42),.acc(r105_42),.res(r105_43),.clk(clk),.wout(w105_43));
	PE pe105_44(.x(x44),.w(w105_43),.acc(r105_43),.res(r105_44),.clk(clk),.wout(w105_44));
	PE pe105_45(.x(x45),.w(w105_44),.acc(r105_44),.res(r105_45),.clk(clk),.wout(w105_45));
	PE pe105_46(.x(x46),.w(w105_45),.acc(r105_45),.res(r105_46),.clk(clk),.wout(w105_46));
	PE pe105_47(.x(x47),.w(w105_46),.acc(r105_46),.res(r105_47),.clk(clk),.wout(w105_47));
	PE pe105_48(.x(x48),.w(w105_47),.acc(r105_47),.res(r105_48),.clk(clk),.wout(w105_48));
	PE pe105_49(.x(x49),.w(w105_48),.acc(r105_48),.res(r105_49),.clk(clk),.wout(w105_49));
	PE pe105_50(.x(x50),.w(w105_49),.acc(r105_49),.res(r105_50),.clk(clk),.wout(w105_50));
	PE pe105_51(.x(x51),.w(w105_50),.acc(r105_50),.res(r105_51),.clk(clk),.wout(w105_51));
	PE pe105_52(.x(x52),.w(w105_51),.acc(r105_51),.res(r105_52),.clk(clk),.wout(w105_52));
	PE pe105_53(.x(x53),.w(w105_52),.acc(r105_52),.res(r105_53),.clk(clk),.wout(w105_53));
	PE pe105_54(.x(x54),.w(w105_53),.acc(r105_53),.res(r105_54),.clk(clk),.wout(w105_54));
	PE pe105_55(.x(x55),.w(w105_54),.acc(r105_54),.res(r105_55),.clk(clk),.wout(w105_55));
	PE pe105_56(.x(x56),.w(w105_55),.acc(r105_55),.res(r105_56),.clk(clk),.wout(w105_56));
	PE pe105_57(.x(x57),.w(w105_56),.acc(r105_56),.res(r105_57),.clk(clk),.wout(w105_57));
	PE pe105_58(.x(x58),.w(w105_57),.acc(r105_57),.res(r105_58),.clk(clk),.wout(w105_58));
	PE pe105_59(.x(x59),.w(w105_58),.acc(r105_58),.res(r105_59),.clk(clk),.wout(w105_59));
	PE pe105_60(.x(x60),.w(w105_59),.acc(r105_59),.res(r105_60),.clk(clk),.wout(w105_60));
	PE pe105_61(.x(x61),.w(w105_60),.acc(r105_60),.res(r105_61),.clk(clk),.wout(w105_61));
	PE pe105_62(.x(x62),.w(w105_61),.acc(r105_61),.res(r105_62),.clk(clk),.wout(w105_62));
	PE pe105_63(.x(x63),.w(w105_62),.acc(r105_62),.res(r105_63),.clk(clk),.wout(w105_63));
	PE pe105_64(.x(x64),.w(w105_63),.acc(r105_63),.res(r105_64),.clk(clk),.wout(w105_64));
	PE pe105_65(.x(x65),.w(w105_64),.acc(r105_64),.res(r105_65),.clk(clk),.wout(w105_65));
	PE pe105_66(.x(x66),.w(w105_65),.acc(r105_65),.res(r105_66),.clk(clk),.wout(w105_66));
	PE pe105_67(.x(x67),.w(w105_66),.acc(r105_66),.res(r105_67),.clk(clk),.wout(w105_67));
	PE pe105_68(.x(x68),.w(w105_67),.acc(r105_67),.res(r105_68),.clk(clk),.wout(w105_68));
	PE pe105_69(.x(x69),.w(w105_68),.acc(r105_68),.res(r105_69),.clk(clk),.wout(w105_69));
	PE pe105_70(.x(x70),.w(w105_69),.acc(r105_69),.res(r105_70),.clk(clk),.wout(w105_70));
	PE pe105_71(.x(x71),.w(w105_70),.acc(r105_70),.res(r105_71),.clk(clk),.wout(w105_71));
	PE pe105_72(.x(x72),.w(w105_71),.acc(r105_71),.res(r105_72),.clk(clk),.wout(w105_72));
	PE pe105_73(.x(x73),.w(w105_72),.acc(r105_72),.res(r105_73),.clk(clk),.wout(w105_73));
	PE pe105_74(.x(x74),.w(w105_73),.acc(r105_73),.res(r105_74),.clk(clk),.wout(w105_74));
	PE pe105_75(.x(x75),.w(w105_74),.acc(r105_74),.res(r105_75),.clk(clk),.wout(w105_75));
	PE pe105_76(.x(x76),.w(w105_75),.acc(r105_75),.res(r105_76),.clk(clk),.wout(w105_76));
	PE pe105_77(.x(x77),.w(w105_76),.acc(r105_76),.res(r105_77),.clk(clk),.wout(w105_77));
	PE pe105_78(.x(x78),.w(w105_77),.acc(r105_77),.res(r105_78),.clk(clk),.wout(w105_78));
	PE pe105_79(.x(x79),.w(w105_78),.acc(r105_78),.res(r105_79),.clk(clk),.wout(w105_79));
	PE pe105_80(.x(x80),.w(w105_79),.acc(r105_79),.res(r105_80),.clk(clk),.wout(w105_80));
	PE pe105_81(.x(x81),.w(w105_80),.acc(r105_80),.res(r105_81),.clk(clk),.wout(w105_81));
	PE pe105_82(.x(x82),.w(w105_81),.acc(r105_81),.res(r105_82),.clk(clk),.wout(w105_82));
	PE pe105_83(.x(x83),.w(w105_82),.acc(r105_82),.res(r105_83),.clk(clk),.wout(w105_83));
	PE pe105_84(.x(x84),.w(w105_83),.acc(r105_83),.res(r105_84),.clk(clk),.wout(w105_84));
	PE pe105_85(.x(x85),.w(w105_84),.acc(r105_84),.res(r105_85),.clk(clk),.wout(w105_85));
	PE pe105_86(.x(x86),.w(w105_85),.acc(r105_85),.res(r105_86),.clk(clk),.wout(w105_86));
	PE pe105_87(.x(x87),.w(w105_86),.acc(r105_86),.res(r105_87),.clk(clk),.wout(w105_87));
	PE pe105_88(.x(x88),.w(w105_87),.acc(r105_87),.res(r105_88),.clk(clk),.wout(w105_88));
	PE pe105_89(.x(x89),.w(w105_88),.acc(r105_88),.res(r105_89),.clk(clk),.wout(w105_89));
	PE pe105_90(.x(x90),.w(w105_89),.acc(r105_89),.res(r105_90),.clk(clk),.wout(w105_90));
	PE pe105_91(.x(x91),.w(w105_90),.acc(r105_90),.res(r105_91),.clk(clk),.wout(w105_91));
	PE pe105_92(.x(x92),.w(w105_91),.acc(r105_91),.res(r105_92),.clk(clk),.wout(w105_92));
	PE pe105_93(.x(x93),.w(w105_92),.acc(r105_92),.res(r105_93),.clk(clk),.wout(w105_93));
	PE pe105_94(.x(x94),.w(w105_93),.acc(r105_93),.res(r105_94),.clk(clk),.wout(w105_94));
	PE pe105_95(.x(x95),.w(w105_94),.acc(r105_94),.res(r105_95),.clk(clk),.wout(w105_95));
	PE pe105_96(.x(x96),.w(w105_95),.acc(r105_95),.res(r105_96),.clk(clk),.wout(w105_96));
	PE pe105_97(.x(x97),.w(w105_96),.acc(r105_96),.res(r105_97),.clk(clk),.wout(w105_97));
	PE pe105_98(.x(x98),.w(w105_97),.acc(r105_97),.res(r105_98),.clk(clk),.wout(w105_98));
	PE pe105_99(.x(x99),.w(w105_98),.acc(r105_98),.res(r105_99),.clk(clk),.wout(w105_99));
	PE pe105_100(.x(x100),.w(w105_99),.acc(r105_99),.res(r105_100),.clk(clk),.wout(w105_100));
	PE pe105_101(.x(x101),.w(w105_100),.acc(r105_100),.res(r105_101),.clk(clk),.wout(w105_101));
	PE pe105_102(.x(x102),.w(w105_101),.acc(r105_101),.res(r105_102),.clk(clk),.wout(w105_102));
	PE pe105_103(.x(x103),.w(w105_102),.acc(r105_102),.res(r105_103),.clk(clk),.wout(w105_103));
	PE pe105_104(.x(x104),.w(w105_103),.acc(r105_103),.res(r105_104),.clk(clk),.wout(w105_104));
	PE pe105_105(.x(x105),.w(w105_104),.acc(r105_104),.res(r105_105),.clk(clk),.wout(w105_105));
	PE pe105_106(.x(x106),.w(w105_105),.acc(r105_105),.res(r105_106),.clk(clk),.wout(w105_106));
	PE pe105_107(.x(x107),.w(w105_106),.acc(r105_106),.res(r105_107),.clk(clk),.wout(w105_107));
	PE pe105_108(.x(x108),.w(w105_107),.acc(r105_107),.res(r105_108),.clk(clk),.wout(w105_108));
	PE pe105_109(.x(x109),.w(w105_108),.acc(r105_108),.res(r105_109),.clk(clk),.wout(w105_109));
	PE pe105_110(.x(x110),.w(w105_109),.acc(r105_109),.res(r105_110),.clk(clk),.wout(w105_110));
	PE pe105_111(.x(x111),.w(w105_110),.acc(r105_110),.res(r105_111),.clk(clk),.wout(w105_111));
	PE pe105_112(.x(x112),.w(w105_111),.acc(r105_111),.res(r105_112),.clk(clk),.wout(w105_112));
	PE pe105_113(.x(x113),.w(w105_112),.acc(r105_112),.res(r105_113),.clk(clk),.wout(w105_113));
	PE pe105_114(.x(x114),.w(w105_113),.acc(r105_113),.res(r105_114),.clk(clk),.wout(w105_114));
	PE pe105_115(.x(x115),.w(w105_114),.acc(r105_114),.res(r105_115),.clk(clk),.wout(w105_115));
	PE pe105_116(.x(x116),.w(w105_115),.acc(r105_115),.res(r105_116),.clk(clk),.wout(w105_116));
	PE pe105_117(.x(x117),.w(w105_116),.acc(r105_116),.res(r105_117),.clk(clk),.wout(w105_117));
	PE pe105_118(.x(x118),.w(w105_117),.acc(r105_117),.res(r105_118),.clk(clk),.wout(w105_118));
	PE pe105_119(.x(x119),.w(w105_118),.acc(r105_118),.res(r105_119),.clk(clk),.wout(w105_119));
	PE pe105_120(.x(x120),.w(w105_119),.acc(r105_119),.res(r105_120),.clk(clk),.wout(w105_120));
	PE pe105_121(.x(x121),.w(w105_120),.acc(r105_120),.res(r105_121),.clk(clk),.wout(w105_121));
	PE pe105_122(.x(x122),.w(w105_121),.acc(r105_121),.res(r105_122),.clk(clk),.wout(w105_122));
	PE pe105_123(.x(x123),.w(w105_122),.acc(r105_122),.res(r105_123),.clk(clk),.wout(w105_123));
	PE pe105_124(.x(x124),.w(w105_123),.acc(r105_123),.res(r105_124),.clk(clk),.wout(w105_124));
	PE pe105_125(.x(x125),.w(w105_124),.acc(r105_124),.res(r105_125),.clk(clk),.wout(w105_125));
	PE pe105_126(.x(x126),.w(w105_125),.acc(r105_125),.res(r105_126),.clk(clk),.wout(w105_126));
	PE pe105_127(.x(x127),.w(w105_126),.acc(r105_126),.res(result105),.clk(clk),.wout(weight105));

	PE pe106_0(.x(x0),.w(w106),.acc(32'h0),.res(r106_0),.clk(clk),.wout(w106_0));
	PE pe106_1(.x(x1),.w(w106_0),.acc(r106_0),.res(r106_1),.clk(clk),.wout(w106_1));
	PE pe106_2(.x(x2),.w(w106_1),.acc(r106_1),.res(r106_2),.clk(clk),.wout(w106_2));
	PE pe106_3(.x(x3),.w(w106_2),.acc(r106_2),.res(r106_3),.clk(clk),.wout(w106_3));
	PE pe106_4(.x(x4),.w(w106_3),.acc(r106_3),.res(r106_4),.clk(clk),.wout(w106_4));
	PE pe106_5(.x(x5),.w(w106_4),.acc(r106_4),.res(r106_5),.clk(clk),.wout(w106_5));
	PE pe106_6(.x(x6),.w(w106_5),.acc(r106_5),.res(r106_6),.clk(clk),.wout(w106_6));
	PE pe106_7(.x(x7),.w(w106_6),.acc(r106_6),.res(r106_7),.clk(clk),.wout(w106_7));
	PE pe106_8(.x(x8),.w(w106_7),.acc(r106_7),.res(r106_8),.clk(clk),.wout(w106_8));
	PE pe106_9(.x(x9),.w(w106_8),.acc(r106_8),.res(r106_9),.clk(clk),.wout(w106_9));
	PE pe106_10(.x(x10),.w(w106_9),.acc(r106_9),.res(r106_10),.clk(clk),.wout(w106_10));
	PE pe106_11(.x(x11),.w(w106_10),.acc(r106_10),.res(r106_11),.clk(clk),.wout(w106_11));
	PE pe106_12(.x(x12),.w(w106_11),.acc(r106_11),.res(r106_12),.clk(clk),.wout(w106_12));
	PE pe106_13(.x(x13),.w(w106_12),.acc(r106_12),.res(r106_13),.clk(clk),.wout(w106_13));
	PE pe106_14(.x(x14),.w(w106_13),.acc(r106_13),.res(r106_14),.clk(clk),.wout(w106_14));
	PE pe106_15(.x(x15),.w(w106_14),.acc(r106_14),.res(r106_15),.clk(clk),.wout(w106_15));
	PE pe106_16(.x(x16),.w(w106_15),.acc(r106_15),.res(r106_16),.clk(clk),.wout(w106_16));
	PE pe106_17(.x(x17),.w(w106_16),.acc(r106_16),.res(r106_17),.clk(clk),.wout(w106_17));
	PE pe106_18(.x(x18),.w(w106_17),.acc(r106_17),.res(r106_18),.clk(clk),.wout(w106_18));
	PE pe106_19(.x(x19),.w(w106_18),.acc(r106_18),.res(r106_19),.clk(clk),.wout(w106_19));
	PE pe106_20(.x(x20),.w(w106_19),.acc(r106_19),.res(r106_20),.clk(clk),.wout(w106_20));
	PE pe106_21(.x(x21),.w(w106_20),.acc(r106_20),.res(r106_21),.clk(clk),.wout(w106_21));
	PE pe106_22(.x(x22),.w(w106_21),.acc(r106_21),.res(r106_22),.clk(clk),.wout(w106_22));
	PE pe106_23(.x(x23),.w(w106_22),.acc(r106_22),.res(r106_23),.clk(clk),.wout(w106_23));
	PE pe106_24(.x(x24),.w(w106_23),.acc(r106_23),.res(r106_24),.clk(clk),.wout(w106_24));
	PE pe106_25(.x(x25),.w(w106_24),.acc(r106_24),.res(r106_25),.clk(clk),.wout(w106_25));
	PE pe106_26(.x(x26),.w(w106_25),.acc(r106_25),.res(r106_26),.clk(clk),.wout(w106_26));
	PE pe106_27(.x(x27),.w(w106_26),.acc(r106_26),.res(r106_27),.clk(clk),.wout(w106_27));
	PE pe106_28(.x(x28),.w(w106_27),.acc(r106_27),.res(r106_28),.clk(clk),.wout(w106_28));
	PE pe106_29(.x(x29),.w(w106_28),.acc(r106_28),.res(r106_29),.clk(clk),.wout(w106_29));
	PE pe106_30(.x(x30),.w(w106_29),.acc(r106_29),.res(r106_30),.clk(clk),.wout(w106_30));
	PE pe106_31(.x(x31),.w(w106_30),.acc(r106_30),.res(r106_31),.clk(clk),.wout(w106_31));
	PE pe106_32(.x(x32),.w(w106_31),.acc(r106_31),.res(r106_32),.clk(clk),.wout(w106_32));
	PE pe106_33(.x(x33),.w(w106_32),.acc(r106_32),.res(r106_33),.clk(clk),.wout(w106_33));
	PE pe106_34(.x(x34),.w(w106_33),.acc(r106_33),.res(r106_34),.clk(clk),.wout(w106_34));
	PE pe106_35(.x(x35),.w(w106_34),.acc(r106_34),.res(r106_35),.clk(clk),.wout(w106_35));
	PE pe106_36(.x(x36),.w(w106_35),.acc(r106_35),.res(r106_36),.clk(clk),.wout(w106_36));
	PE pe106_37(.x(x37),.w(w106_36),.acc(r106_36),.res(r106_37),.clk(clk),.wout(w106_37));
	PE pe106_38(.x(x38),.w(w106_37),.acc(r106_37),.res(r106_38),.clk(clk),.wout(w106_38));
	PE pe106_39(.x(x39),.w(w106_38),.acc(r106_38),.res(r106_39),.clk(clk),.wout(w106_39));
	PE pe106_40(.x(x40),.w(w106_39),.acc(r106_39),.res(r106_40),.clk(clk),.wout(w106_40));
	PE pe106_41(.x(x41),.w(w106_40),.acc(r106_40),.res(r106_41),.clk(clk),.wout(w106_41));
	PE pe106_42(.x(x42),.w(w106_41),.acc(r106_41),.res(r106_42),.clk(clk),.wout(w106_42));
	PE pe106_43(.x(x43),.w(w106_42),.acc(r106_42),.res(r106_43),.clk(clk),.wout(w106_43));
	PE pe106_44(.x(x44),.w(w106_43),.acc(r106_43),.res(r106_44),.clk(clk),.wout(w106_44));
	PE pe106_45(.x(x45),.w(w106_44),.acc(r106_44),.res(r106_45),.clk(clk),.wout(w106_45));
	PE pe106_46(.x(x46),.w(w106_45),.acc(r106_45),.res(r106_46),.clk(clk),.wout(w106_46));
	PE pe106_47(.x(x47),.w(w106_46),.acc(r106_46),.res(r106_47),.clk(clk),.wout(w106_47));
	PE pe106_48(.x(x48),.w(w106_47),.acc(r106_47),.res(r106_48),.clk(clk),.wout(w106_48));
	PE pe106_49(.x(x49),.w(w106_48),.acc(r106_48),.res(r106_49),.clk(clk),.wout(w106_49));
	PE pe106_50(.x(x50),.w(w106_49),.acc(r106_49),.res(r106_50),.clk(clk),.wout(w106_50));
	PE pe106_51(.x(x51),.w(w106_50),.acc(r106_50),.res(r106_51),.clk(clk),.wout(w106_51));
	PE pe106_52(.x(x52),.w(w106_51),.acc(r106_51),.res(r106_52),.clk(clk),.wout(w106_52));
	PE pe106_53(.x(x53),.w(w106_52),.acc(r106_52),.res(r106_53),.clk(clk),.wout(w106_53));
	PE pe106_54(.x(x54),.w(w106_53),.acc(r106_53),.res(r106_54),.clk(clk),.wout(w106_54));
	PE pe106_55(.x(x55),.w(w106_54),.acc(r106_54),.res(r106_55),.clk(clk),.wout(w106_55));
	PE pe106_56(.x(x56),.w(w106_55),.acc(r106_55),.res(r106_56),.clk(clk),.wout(w106_56));
	PE pe106_57(.x(x57),.w(w106_56),.acc(r106_56),.res(r106_57),.clk(clk),.wout(w106_57));
	PE pe106_58(.x(x58),.w(w106_57),.acc(r106_57),.res(r106_58),.clk(clk),.wout(w106_58));
	PE pe106_59(.x(x59),.w(w106_58),.acc(r106_58),.res(r106_59),.clk(clk),.wout(w106_59));
	PE pe106_60(.x(x60),.w(w106_59),.acc(r106_59),.res(r106_60),.clk(clk),.wout(w106_60));
	PE pe106_61(.x(x61),.w(w106_60),.acc(r106_60),.res(r106_61),.clk(clk),.wout(w106_61));
	PE pe106_62(.x(x62),.w(w106_61),.acc(r106_61),.res(r106_62),.clk(clk),.wout(w106_62));
	PE pe106_63(.x(x63),.w(w106_62),.acc(r106_62),.res(r106_63),.clk(clk),.wout(w106_63));
	PE pe106_64(.x(x64),.w(w106_63),.acc(r106_63),.res(r106_64),.clk(clk),.wout(w106_64));
	PE pe106_65(.x(x65),.w(w106_64),.acc(r106_64),.res(r106_65),.clk(clk),.wout(w106_65));
	PE pe106_66(.x(x66),.w(w106_65),.acc(r106_65),.res(r106_66),.clk(clk),.wout(w106_66));
	PE pe106_67(.x(x67),.w(w106_66),.acc(r106_66),.res(r106_67),.clk(clk),.wout(w106_67));
	PE pe106_68(.x(x68),.w(w106_67),.acc(r106_67),.res(r106_68),.clk(clk),.wout(w106_68));
	PE pe106_69(.x(x69),.w(w106_68),.acc(r106_68),.res(r106_69),.clk(clk),.wout(w106_69));
	PE pe106_70(.x(x70),.w(w106_69),.acc(r106_69),.res(r106_70),.clk(clk),.wout(w106_70));
	PE pe106_71(.x(x71),.w(w106_70),.acc(r106_70),.res(r106_71),.clk(clk),.wout(w106_71));
	PE pe106_72(.x(x72),.w(w106_71),.acc(r106_71),.res(r106_72),.clk(clk),.wout(w106_72));
	PE pe106_73(.x(x73),.w(w106_72),.acc(r106_72),.res(r106_73),.clk(clk),.wout(w106_73));
	PE pe106_74(.x(x74),.w(w106_73),.acc(r106_73),.res(r106_74),.clk(clk),.wout(w106_74));
	PE pe106_75(.x(x75),.w(w106_74),.acc(r106_74),.res(r106_75),.clk(clk),.wout(w106_75));
	PE pe106_76(.x(x76),.w(w106_75),.acc(r106_75),.res(r106_76),.clk(clk),.wout(w106_76));
	PE pe106_77(.x(x77),.w(w106_76),.acc(r106_76),.res(r106_77),.clk(clk),.wout(w106_77));
	PE pe106_78(.x(x78),.w(w106_77),.acc(r106_77),.res(r106_78),.clk(clk),.wout(w106_78));
	PE pe106_79(.x(x79),.w(w106_78),.acc(r106_78),.res(r106_79),.clk(clk),.wout(w106_79));
	PE pe106_80(.x(x80),.w(w106_79),.acc(r106_79),.res(r106_80),.clk(clk),.wout(w106_80));
	PE pe106_81(.x(x81),.w(w106_80),.acc(r106_80),.res(r106_81),.clk(clk),.wout(w106_81));
	PE pe106_82(.x(x82),.w(w106_81),.acc(r106_81),.res(r106_82),.clk(clk),.wout(w106_82));
	PE pe106_83(.x(x83),.w(w106_82),.acc(r106_82),.res(r106_83),.clk(clk),.wout(w106_83));
	PE pe106_84(.x(x84),.w(w106_83),.acc(r106_83),.res(r106_84),.clk(clk),.wout(w106_84));
	PE pe106_85(.x(x85),.w(w106_84),.acc(r106_84),.res(r106_85),.clk(clk),.wout(w106_85));
	PE pe106_86(.x(x86),.w(w106_85),.acc(r106_85),.res(r106_86),.clk(clk),.wout(w106_86));
	PE pe106_87(.x(x87),.w(w106_86),.acc(r106_86),.res(r106_87),.clk(clk),.wout(w106_87));
	PE pe106_88(.x(x88),.w(w106_87),.acc(r106_87),.res(r106_88),.clk(clk),.wout(w106_88));
	PE pe106_89(.x(x89),.w(w106_88),.acc(r106_88),.res(r106_89),.clk(clk),.wout(w106_89));
	PE pe106_90(.x(x90),.w(w106_89),.acc(r106_89),.res(r106_90),.clk(clk),.wout(w106_90));
	PE pe106_91(.x(x91),.w(w106_90),.acc(r106_90),.res(r106_91),.clk(clk),.wout(w106_91));
	PE pe106_92(.x(x92),.w(w106_91),.acc(r106_91),.res(r106_92),.clk(clk),.wout(w106_92));
	PE pe106_93(.x(x93),.w(w106_92),.acc(r106_92),.res(r106_93),.clk(clk),.wout(w106_93));
	PE pe106_94(.x(x94),.w(w106_93),.acc(r106_93),.res(r106_94),.clk(clk),.wout(w106_94));
	PE pe106_95(.x(x95),.w(w106_94),.acc(r106_94),.res(r106_95),.clk(clk),.wout(w106_95));
	PE pe106_96(.x(x96),.w(w106_95),.acc(r106_95),.res(r106_96),.clk(clk),.wout(w106_96));
	PE pe106_97(.x(x97),.w(w106_96),.acc(r106_96),.res(r106_97),.clk(clk),.wout(w106_97));
	PE pe106_98(.x(x98),.w(w106_97),.acc(r106_97),.res(r106_98),.clk(clk),.wout(w106_98));
	PE pe106_99(.x(x99),.w(w106_98),.acc(r106_98),.res(r106_99),.clk(clk),.wout(w106_99));
	PE pe106_100(.x(x100),.w(w106_99),.acc(r106_99),.res(r106_100),.clk(clk),.wout(w106_100));
	PE pe106_101(.x(x101),.w(w106_100),.acc(r106_100),.res(r106_101),.clk(clk),.wout(w106_101));
	PE pe106_102(.x(x102),.w(w106_101),.acc(r106_101),.res(r106_102),.clk(clk),.wout(w106_102));
	PE pe106_103(.x(x103),.w(w106_102),.acc(r106_102),.res(r106_103),.clk(clk),.wout(w106_103));
	PE pe106_104(.x(x104),.w(w106_103),.acc(r106_103),.res(r106_104),.clk(clk),.wout(w106_104));
	PE pe106_105(.x(x105),.w(w106_104),.acc(r106_104),.res(r106_105),.clk(clk),.wout(w106_105));
	PE pe106_106(.x(x106),.w(w106_105),.acc(r106_105),.res(r106_106),.clk(clk),.wout(w106_106));
	PE pe106_107(.x(x107),.w(w106_106),.acc(r106_106),.res(r106_107),.clk(clk),.wout(w106_107));
	PE pe106_108(.x(x108),.w(w106_107),.acc(r106_107),.res(r106_108),.clk(clk),.wout(w106_108));
	PE pe106_109(.x(x109),.w(w106_108),.acc(r106_108),.res(r106_109),.clk(clk),.wout(w106_109));
	PE pe106_110(.x(x110),.w(w106_109),.acc(r106_109),.res(r106_110),.clk(clk),.wout(w106_110));
	PE pe106_111(.x(x111),.w(w106_110),.acc(r106_110),.res(r106_111),.clk(clk),.wout(w106_111));
	PE pe106_112(.x(x112),.w(w106_111),.acc(r106_111),.res(r106_112),.clk(clk),.wout(w106_112));
	PE pe106_113(.x(x113),.w(w106_112),.acc(r106_112),.res(r106_113),.clk(clk),.wout(w106_113));
	PE pe106_114(.x(x114),.w(w106_113),.acc(r106_113),.res(r106_114),.clk(clk),.wout(w106_114));
	PE pe106_115(.x(x115),.w(w106_114),.acc(r106_114),.res(r106_115),.clk(clk),.wout(w106_115));
	PE pe106_116(.x(x116),.w(w106_115),.acc(r106_115),.res(r106_116),.clk(clk),.wout(w106_116));
	PE pe106_117(.x(x117),.w(w106_116),.acc(r106_116),.res(r106_117),.clk(clk),.wout(w106_117));
	PE pe106_118(.x(x118),.w(w106_117),.acc(r106_117),.res(r106_118),.clk(clk),.wout(w106_118));
	PE pe106_119(.x(x119),.w(w106_118),.acc(r106_118),.res(r106_119),.clk(clk),.wout(w106_119));
	PE pe106_120(.x(x120),.w(w106_119),.acc(r106_119),.res(r106_120),.clk(clk),.wout(w106_120));
	PE pe106_121(.x(x121),.w(w106_120),.acc(r106_120),.res(r106_121),.clk(clk),.wout(w106_121));
	PE pe106_122(.x(x122),.w(w106_121),.acc(r106_121),.res(r106_122),.clk(clk),.wout(w106_122));
	PE pe106_123(.x(x123),.w(w106_122),.acc(r106_122),.res(r106_123),.clk(clk),.wout(w106_123));
	PE pe106_124(.x(x124),.w(w106_123),.acc(r106_123),.res(r106_124),.clk(clk),.wout(w106_124));
	PE pe106_125(.x(x125),.w(w106_124),.acc(r106_124),.res(r106_125),.clk(clk),.wout(w106_125));
	PE pe106_126(.x(x126),.w(w106_125),.acc(r106_125),.res(r106_126),.clk(clk),.wout(w106_126));
	PE pe106_127(.x(x127),.w(w106_126),.acc(r106_126),.res(result106),.clk(clk),.wout(weight106));

	PE pe107_0(.x(x0),.w(w107),.acc(32'h0),.res(r107_0),.clk(clk),.wout(w107_0));
	PE pe107_1(.x(x1),.w(w107_0),.acc(r107_0),.res(r107_1),.clk(clk),.wout(w107_1));
	PE pe107_2(.x(x2),.w(w107_1),.acc(r107_1),.res(r107_2),.clk(clk),.wout(w107_2));
	PE pe107_3(.x(x3),.w(w107_2),.acc(r107_2),.res(r107_3),.clk(clk),.wout(w107_3));
	PE pe107_4(.x(x4),.w(w107_3),.acc(r107_3),.res(r107_4),.clk(clk),.wout(w107_4));
	PE pe107_5(.x(x5),.w(w107_4),.acc(r107_4),.res(r107_5),.clk(clk),.wout(w107_5));
	PE pe107_6(.x(x6),.w(w107_5),.acc(r107_5),.res(r107_6),.clk(clk),.wout(w107_6));
	PE pe107_7(.x(x7),.w(w107_6),.acc(r107_6),.res(r107_7),.clk(clk),.wout(w107_7));
	PE pe107_8(.x(x8),.w(w107_7),.acc(r107_7),.res(r107_8),.clk(clk),.wout(w107_8));
	PE pe107_9(.x(x9),.w(w107_8),.acc(r107_8),.res(r107_9),.clk(clk),.wout(w107_9));
	PE pe107_10(.x(x10),.w(w107_9),.acc(r107_9),.res(r107_10),.clk(clk),.wout(w107_10));
	PE pe107_11(.x(x11),.w(w107_10),.acc(r107_10),.res(r107_11),.clk(clk),.wout(w107_11));
	PE pe107_12(.x(x12),.w(w107_11),.acc(r107_11),.res(r107_12),.clk(clk),.wout(w107_12));
	PE pe107_13(.x(x13),.w(w107_12),.acc(r107_12),.res(r107_13),.clk(clk),.wout(w107_13));
	PE pe107_14(.x(x14),.w(w107_13),.acc(r107_13),.res(r107_14),.clk(clk),.wout(w107_14));
	PE pe107_15(.x(x15),.w(w107_14),.acc(r107_14),.res(r107_15),.clk(clk),.wout(w107_15));
	PE pe107_16(.x(x16),.w(w107_15),.acc(r107_15),.res(r107_16),.clk(clk),.wout(w107_16));
	PE pe107_17(.x(x17),.w(w107_16),.acc(r107_16),.res(r107_17),.clk(clk),.wout(w107_17));
	PE pe107_18(.x(x18),.w(w107_17),.acc(r107_17),.res(r107_18),.clk(clk),.wout(w107_18));
	PE pe107_19(.x(x19),.w(w107_18),.acc(r107_18),.res(r107_19),.clk(clk),.wout(w107_19));
	PE pe107_20(.x(x20),.w(w107_19),.acc(r107_19),.res(r107_20),.clk(clk),.wout(w107_20));
	PE pe107_21(.x(x21),.w(w107_20),.acc(r107_20),.res(r107_21),.clk(clk),.wout(w107_21));
	PE pe107_22(.x(x22),.w(w107_21),.acc(r107_21),.res(r107_22),.clk(clk),.wout(w107_22));
	PE pe107_23(.x(x23),.w(w107_22),.acc(r107_22),.res(r107_23),.clk(clk),.wout(w107_23));
	PE pe107_24(.x(x24),.w(w107_23),.acc(r107_23),.res(r107_24),.clk(clk),.wout(w107_24));
	PE pe107_25(.x(x25),.w(w107_24),.acc(r107_24),.res(r107_25),.clk(clk),.wout(w107_25));
	PE pe107_26(.x(x26),.w(w107_25),.acc(r107_25),.res(r107_26),.clk(clk),.wout(w107_26));
	PE pe107_27(.x(x27),.w(w107_26),.acc(r107_26),.res(r107_27),.clk(clk),.wout(w107_27));
	PE pe107_28(.x(x28),.w(w107_27),.acc(r107_27),.res(r107_28),.clk(clk),.wout(w107_28));
	PE pe107_29(.x(x29),.w(w107_28),.acc(r107_28),.res(r107_29),.clk(clk),.wout(w107_29));
	PE pe107_30(.x(x30),.w(w107_29),.acc(r107_29),.res(r107_30),.clk(clk),.wout(w107_30));
	PE pe107_31(.x(x31),.w(w107_30),.acc(r107_30),.res(r107_31),.clk(clk),.wout(w107_31));
	PE pe107_32(.x(x32),.w(w107_31),.acc(r107_31),.res(r107_32),.clk(clk),.wout(w107_32));
	PE pe107_33(.x(x33),.w(w107_32),.acc(r107_32),.res(r107_33),.clk(clk),.wout(w107_33));
	PE pe107_34(.x(x34),.w(w107_33),.acc(r107_33),.res(r107_34),.clk(clk),.wout(w107_34));
	PE pe107_35(.x(x35),.w(w107_34),.acc(r107_34),.res(r107_35),.clk(clk),.wout(w107_35));
	PE pe107_36(.x(x36),.w(w107_35),.acc(r107_35),.res(r107_36),.clk(clk),.wout(w107_36));
	PE pe107_37(.x(x37),.w(w107_36),.acc(r107_36),.res(r107_37),.clk(clk),.wout(w107_37));
	PE pe107_38(.x(x38),.w(w107_37),.acc(r107_37),.res(r107_38),.clk(clk),.wout(w107_38));
	PE pe107_39(.x(x39),.w(w107_38),.acc(r107_38),.res(r107_39),.clk(clk),.wout(w107_39));
	PE pe107_40(.x(x40),.w(w107_39),.acc(r107_39),.res(r107_40),.clk(clk),.wout(w107_40));
	PE pe107_41(.x(x41),.w(w107_40),.acc(r107_40),.res(r107_41),.clk(clk),.wout(w107_41));
	PE pe107_42(.x(x42),.w(w107_41),.acc(r107_41),.res(r107_42),.clk(clk),.wout(w107_42));
	PE pe107_43(.x(x43),.w(w107_42),.acc(r107_42),.res(r107_43),.clk(clk),.wout(w107_43));
	PE pe107_44(.x(x44),.w(w107_43),.acc(r107_43),.res(r107_44),.clk(clk),.wout(w107_44));
	PE pe107_45(.x(x45),.w(w107_44),.acc(r107_44),.res(r107_45),.clk(clk),.wout(w107_45));
	PE pe107_46(.x(x46),.w(w107_45),.acc(r107_45),.res(r107_46),.clk(clk),.wout(w107_46));
	PE pe107_47(.x(x47),.w(w107_46),.acc(r107_46),.res(r107_47),.clk(clk),.wout(w107_47));
	PE pe107_48(.x(x48),.w(w107_47),.acc(r107_47),.res(r107_48),.clk(clk),.wout(w107_48));
	PE pe107_49(.x(x49),.w(w107_48),.acc(r107_48),.res(r107_49),.clk(clk),.wout(w107_49));
	PE pe107_50(.x(x50),.w(w107_49),.acc(r107_49),.res(r107_50),.clk(clk),.wout(w107_50));
	PE pe107_51(.x(x51),.w(w107_50),.acc(r107_50),.res(r107_51),.clk(clk),.wout(w107_51));
	PE pe107_52(.x(x52),.w(w107_51),.acc(r107_51),.res(r107_52),.clk(clk),.wout(w107_52));
	PE pe107_53(.x(x53),.w(w107_52),.acc(r107_52),.res(r107_53),.clk(clk),.wout(w107_53));
	PE pe107_54(.x(x54),.w(w107_53),.acc(r107_53),.res(r107_54),.clk(clk),.wout(w107_54));
	PE pe107_55(.x(x55),.w(w107_54),.acc(r107_54),.res(r107_55),.clk(clk),.wout(w107_55));
	PE pe107_56(.x(x56),.w(w107_55),.acc(r107_55),.res(r107_56),.clk(clk),.wout(w107_56));
	PE pe107_57(.x(x57),.w(w107_56),.acc(r107_56),.res(r107_57),.clk(clk),.wout(w107_57));
	PE pe107_58(.x(x58),.w(w107_57),.acc(r107_57),.res(r107_58),.clk(clk),.wout(w107_58));
	PE pe107_59(.x(x59),.w(w107_58),.acc(r107_58),.res(r107_59),.clk(clk),.wout(w107_59));
	PE pe107_60(.x(x60),.w(w107_59),.acc(r107_59),.res(r107_60),.clk(clk),.wout(w107_60));
	PE pe107_61(.x(x61),.w(w107_60),.acc(r107_60),.res(r107_61),.clk(clk),.wout(w107_61));
	PE pe107_62(.x(x62),.w(w107_61),.acc(r107_61),.res(r107_62),.clk(clk),.wout(w107_62));
	PE pe107_63(.x(x63),.w(w107_62),.acc(r107_62),.res(r107_63),.clk(clk),.wout(w107_63));
	PE pe107_64(.x(x64),.w(w107_63),.acc(r107_63),.res(r107_64),.clk(clk),.wout(w107_64));
	PE pe107_65(.x(x65),.w(w107_64),.acc(r107_64),.res(r107_65),.clk(clk),.wout(w107_65));
	PE pe107_66(.x(x66),.w(w107_65),.acc(r107_65),.res(r107_66),.clk(clk),.wout(w107_66));
	PE pe107_67(.x(x67),.w(w107_66),.acc(r107_66),.res(r107_67),.clk(clk),.wout(w107_67));
	PE pe107_68(.x(x68),.w(w107_67),.acc(r107_67),.res(r107_68),.clk(clk),.wout(w107_68));
	PE pe107_69(.x(x69),.w(w107_68),.acc(r107_68),.res(r107_69),.clk(clk),.wout(w107_69));
	PE pe107_70(.x(x70),.w(w107_69),.acc(r107_69),.res(r107_70),.clk(clk),.wout(w107_70));
	PE pe107_71(.x(x71),.w(w107_70),.acc(r107_70),.res(r107_71),.clk(clk),.wout(w107_71));
	PE pe107_72(.x(x72),.w(w107_71),.acc(r107_71),.res(r107_72),.clk(clk),.wout(w107_72));
	PE pe107_73(.x(x73),.w(w107_72),.acc(r107_72),.res(r107_73),.clk(clk),.wout(w107_73));
	PE pe107_74(.x(x74),.w(w107_73),.acc(r107_73),.res(r107_74),.clk(clk),.wout(w107_74));
	PE pe107_75(.x(x75),.w(w107_74),.acc(r107_74),.res(r107_75),.clk(clk),.wout(w107_75));
	PE pe107_76(.x(x76),.w(w107_75),.acc(r107_75),.res(r107_76),.clk(clk),.wout(w107_76));
	PE pe107_77(.x(x77),.w(w107_76),.acc(r107_76),.res(r107_77),.clk(clk),.wout(w107_77));
	PE pe107_78(.x(x78),.w(w107_77),.acc(r107_77),.res(r107_78),.clk(clk),.wout(w107_78));
	PE pe107_79(.x(x79),.w(w107_78),.acc(r107_78),.res(r107_79),.clk(clk),.wout(w107_79));
	PE pe107_80(.x(x80),.w(w107_79),.acc(r107_79),.res(r107_80),.clk(clk),.wout(w107_80));
	PE pe107_81(.x(x81),.w(w107_80),.acc(r107_80),.res(r107_81),.clk(clk),.wout(w107_81));
	PE pe107_82(.x(x82),.w(w107_81),.acc(r107_81),.res(r107_82),.clk(clk),.wout(w107_82));
	PE pe107_83(.x(x83),.w(w107_82),.acc(r107_82),.res(r107_83),.clk(clk),.wout(w107_83));
	PE pe107_84(.x(x84),.w(w107_83),.acc(r107_83),.res(r107_84),.clk(clk),.wout(w107_84));
	PE pe107_85(.x(x85),.w(w107_84),.acc(r107_84),.res(r107_85),.clk(clk),.wout(w107_85));
	PE pe107_86(.x(x86),.w(w107_85),.acc(r107_85),.res(r107_86),.clk(clk),.wout(w107_86));
	PE pe107_87(.x(x87),.w(w107_86),.acc(r107_86),.res(r107_87),.clk(clk),.wout(w107_87));
	PE pe107_88(.x(x88),.w(w107_87),.acc(r107_87),.res(r107_88),.clk(clk),.wout(w107_88));
	PE pe107_89(.x(x89),.w(w107_88),.acc(r107_88),.res(r107_89),.clk(clk),.wout(w107_89));
	PE pe107_90(.x(x90),.w(w107_89),.acc(r107_89),.res(r107_90),.clk(clk),.wout(w107_90));
	PE pe107_91(.x(x91),.w(w107_90),.acc(r107_90),.res(r107_91),.clk(clk),.wout(w107_91));
	PE pe107_92(.x(x92),.w(w107_91),.acc(r107_91),.res(r107_92),.clk(clk),.wout(w107_92));
	PE pe107_93(.x(x93),.w(w107_92),.acc(r107_92),.res(r107_93),.clk(clk),.wout(w107_93));
	PE pe107_94(.x(x94),.w(w107_93),.acc(r107_93),.res(r107_94),.clk(clk),.wout(w107_94));
	PE pe107_95(.x(x95),.w(w107_94),.acc(r107_94),.res(r107_95),.clk(clk),.wout(w107_95));
	PE pe107_96(.x(x96),.w(w107_95),.acc(r107_95),.res(r107_96),.clk(clk),.wout(w107_96));
	PE pe107_97(.x(x97),.w(w107_96),.acc(r107_96),.res(r107_97),.clk(clk),.wout(w107_97));
	PE pe107_98(.x(x98),.w(w107_97),.acc(r107_97),.res(r107_98),.clk(clk),.wout(w107_98));
	PE pe107_99(.x(x99),.w(w107_98),.acc(r107_98),.res(r107_99),.clk(clk),.wout(w107_99));
	PE pe107_100(.x(x100),.w(w107_99),.acc(r107_99),.res(r107_100),.clk(clk),.wout(w107_100));
	PE pe107_101(.x(x101),.w(w107_100),.acc(r107_100),.res(r107_101),.clk(clk),.wout(w107_101));
	PE pe107_102(.x(x102),.w(w107_101),.acc(r107_101),.res(r107_102),.clk(clk),.wout(w107_102));
	PE pe107_103(.x(x103),.w(w107_102),.acc(r107_102),.res(r107_103),.clk(clk),.wout(w107_103));
	PE pe107_104(.x(x104),.w(w107_103),.acc(r107_103),.res(r107_104),.clk(clk),.wout(w107_104));
	PE pe107_105(.x(x105),.w(w107_104),.acc(r107_104),.res(r107_105),.clk(clk),.wout(w107_105));
	PE pe107_106(.x(x106),.w(w107_105),.acc(r107_105),.res(r107_106),.clk(clk),.wout(w107_106));
	PE pe107_107(.x(x107),.w(w107_106),.acc(r107_106),.res(r107_107),.clk(clk),.wout(w107_107));
	PE pe107_108(.x(x108),.w(w107_107),.acc(r107_107),.res(r107_108),.clk(clk),.wout(w107_108));
	PE pe107_109(.x(x109),.w(w107_108),.acc(r107_108),.res(r107_109),.clk(clk),.wout(w107_109));
	PE pe107_110(.x(x110),.w(w107_109),.acc(r107_109),.res(r107_110),.clk(clk),.wout(w107_110));
	PE pe107_111(.x(x111),.w(w107_110),.acc(r107_110),.res(r107_111),.clk(clk),.wout(w107_111));
	PE pe107_112(.x(x112),.w(w107_111),.acc(r107_111),.res(r107_112),.clk(clk),.wout(w107_112));
	PE pe107_113(.x(x113),.w(w107_112),.acc(r107_112),.res(r107_113),.clk(clk),.wout(w107_113));
	PE pe107_114(.x(x114),.w(w107_113),.acc(r107_113),.res(r107_114),.clk(clk),.wout(w107_114));
	PE pe107_115(.x(x115),.w(w107_114),.acc(r107_114),.res(r107_115),.clk(clk),.wout(w107_115));
	PE pe107_116(.x(x116),.w(w107_115),.acc(r107_115),.res(r107_116),.clk(clk),.wout(w107_116));
	PE pe107_117(.x(x117),.w(w107_116),.acc(r107_116),.res(r107_117),.clk(clk),.wout(w107_117));
	PE pe107_118(.x(x118),.w(w107_117),.acc(r107_117),.res(r107_118),.clk(clk),.wout(w107_118));
	PE pe107_119(.x(x119),.w(w107_118),.acc(r107_118),.res(r107_119),.clk(clk),.wout(w107_119));
	PE pe107_120(.x(x120),.w(w107_119),.acc(r107_119),.res(r107_120),.clk(clk),.wout(w107_120));
	PE pe107_121(.x(x121),.w(w107_120),.acc(r107_120),.res(r107_121),.clk(clk),.wout(w107_121));
	PE pe107_122(.x(x122),.w(w107_121),.acc(r107_121),.res(r107_122),.clk(clk),.wout(w107_122));
	PE pe107_123(.x(x123),.w(w107_122),.acc(r107_122),.res(r107_123),.clk(clk),.wout(w107_123));
	PE pe107_124(.x(x124),.w(w107_123),.acc(r107_123),.res(r107_124),.clk(clk),.wout(w107_124));
	PE pe107_125(.x(x125),.w(w107_124),.acc(r107_124),.res(r107_125),.clk(clk),.wout(w107_125));
	PE pe107_126(.x(x126),.w(w107_125),.acc(r107_125),.res(r107_126),.clk(clk),.wout(w107_126));
	PE pe107_127(.x(x127),.w(w107_126),.acc(r107_126),.res(result107),.clk(clk),.wout(weight107));

	PE pe108_0(.x(x0),.w(w108),.acc(32'h0),.res(r108_0),.clk(clk),.wout(w108_0));
	PE pe108_1(.x(x1),.w(w108_0),.acc(r108_0),.res(r108_1),.clk(clk),.wout(w108_1));
	PE pe108_2(.x(x2),.w(w108_1),.acc(r108_1),.res(r108_2),.clk(clk),.wout(w108_2));
	PE pe108_3(.x(x3),.w(w108_2),.acc(r108_2),.res(r108_3),.clk(clk),.wout(w108_3));
	PE pe108_4(.x(x4),.w(w108_3),.acc(r108_3),.res(r108_4),.clk(clk),.wout(w108_4));
	PE pe108_5(.x(x5),.w(w108_4),.acc(r108_4),.res(r108_5),.clk(clk),.wout(w108_5));
	PE pe108_6(.x(x6),.w(w108_5),.acc(r108_5),.res(r108_6),.clk(clk),.wout(w108_6));
	PE pe108_7(.x(x7),.w(w108_6),.acc(r108_6),.res(r108_7),.clk(clk),.wout(w108_7));
	PE pe108_8(.x(x8),.w(w108_7),.acc(r108_7),.res(r108_8),.clk(clk),.wout(w108_8));
	PE pe108_9(.x(x9),.w(w108_8),.acc(r108_8),.res(r108_9),.clk(clk),.wout(w108_9));
	PE pe108_10(.x(x10),.w(w108_9),.acc(r108_9),.res(r108_10),.clk(clk),.wout(w108_10));
	PE pe108_11(.x(x11),.w(w108_10),.acc(r108_10),.res(r108_11),.clk(clk),.wout(w108_11));
	PE pe108_12(.x(x12),.w(w108_11),.acc(r108_11),.res(r108_12),.clk(clk),.wout(w108_12));
	PE pe108_13(.x(x13),.w(w108_12),.acc(r108_12),.res(r108_13),.clk(clk),.wout(w108_13));
	PE pe108_14(.x(x14),.w(w108_13),.acc(r108_13),.res(r108_14),.clk(clk),.wout(w108_14));
	PE pe108_15(.x(x15),.w(w108_14),.acc(r108_14),.res(r108_15),.clk(clk),.wout(w108_15));
	PE pe108_16(.x(x16),.w(w108_15),.acc(r108_15),.res(r108_16),.clk(clk),.wout(w108_16));
	PE pe108_17(.x(x17),.w(w108_16),.acc(r108_16),.res(r108_17),.clk(clk),.wout(w108_17));
	PE pe108_18(.x(x18),.w(w108_17),.acc(r108_17),.res(r108_18),.clk(clk),.wout(w108_18));
	PE pe108_19(.x(x19),.w(w108_18),.acc(r108_18),.res(r108_19),.clk(clk),.wout(w108_19));
	PE pe108_20(.x(x20),.w(w108_19),.acc(r108_19),.res(r108_20),.clk(clk),.wout(w108_20));
	PE pe108_21(.x(x21),.w(w108_20),.acc(r108_20),.res(r108_21),.clk(clk),.wout(w108_21));
	PE pe108_22(.x(x22),.w(w108_21),.acc(r108_21),.res(r108_22),.clk(clk),.wout(w108_22));
	PE pe108_23(.x(x23),.w(w108_22),.acc(r108_22),.res(r108_23),.clk(clk),.wout(w108_23));
	PE pe108_24(.x(x24),.w(w108_23),.acc(r108_23),.res(r108_24),.clk(clk),.wout(w108_24));
	PE pe108_25(.x(x25),.w(w108_24),.acc(r108_24),.res(r108_25),.clk(clk),.wout(w108_25));
	PE pe108_26(.x(x26),.w(w108_25),.acc(r108_25),.res(r108_26),.clk(clk),.wout(w108_26));
	PE pe108_27(.x(x27),.w(w108_26),.acc(r108_26),.res(r108_27),.clk(clk),.wout(w108_27));
	PE pe108_28(.x(x28),.w(w108_27),.acc(r108_27),.res(r108_28),.clk(clk),.wout(w108_28));
	PE pe108_29(.x(x29),.w(w108_28),.acc(r108_28),.res(r108_29),.clk(clk),.wout(w108_29));
	PE pe108_30(.x(x30),.w(w108_29),.acc(r108_29),.res(r108_30),.clk(clk),.wout(w108_30));
	PE pe108_31(.x(x31),.w(w108_30),.acc(r108_30),.res(r108_31),.clk(clk),.wout(w108_31));
	PE pe108_32(.x(x32),.w(w108_31),.acc(r108_31),.res(r108_32),.clk(clk),.wout(w108_32));
	PE pe108_33(.x(x33),.w(w108_32),.acc(r108_32),.res(r108_33),.clk(clk),.wout(w108_33));
	PE pe108_34(.x(x34),.w(w108_33),.acc(r108_33),.res(r108_34),.clk(clk),.wout(w108_34));
	PE pe108_35(.x(x35),.w(w108_34),.acc(r108_34),.res(r108_35),.clk(clk),.wout(w108_35));
	PE pe108_36(.x(x36),.w(w108_35),.acc(r108_35),.res(r108_36),.clk(clk),.wout(w108_36));
	PE pe108_37(.x(x37),.w(w108_36),.acc(r108_36),.res(r108_37),.clk(clk),.wout(w108_37));
	PE pe108_38(.x(x38),.w(w108_37),.acc(r108_37),.res(r108_38),.clk(clk),.wout(w108_38));
	PE pe108_39(.x(x39),.w(w108_38),.acc(r108_38),.res(r108_39),.clk(clk),.wout(w108_39));
	PE pe108_40(.x(x40),.w(w108_39),.acc(r108_39),.res(r108_40),.clk(clk),.wout(w108_40));
	PE pe108_41(.x(x41),.w(w108_40),.acc(r108_40),.res(r108_41),.clk(clk),.wout(w108_41));
	PE pe108_42(.x(x42),.w(w108_41),.acc(r108_41),.res(r108_42),.clk(clk),.wout(w108_42));
	PE pe108_43(.x(x43),.w(w108_42),.acc(r108_42),.res(r108_43),.clk(clk),.wout(w108_43));
	PE pe108_44(.x(x44),.w(w108_43),.acc(r108_43),.res(r108_44),.clk(clk),.wout(w108_44));
	PE pe108_45(.x(x45),.w(w108_44),.acc(r108_44),.res(r108_45),.clk(clk),.wout(w108_45));
	PE pe108_46(.x(x46),.w(w108_45),.acc(r108_45),.res(r108_46),.clk(clk),.wout(w108_46));
	PE pe108_47(.x(x47),.w(w108_46),.acc(r108_46),.res(r108_47),.clk(clk),.wout(w108_47));
	PE pe108_48(.x(x48),.w(w108_47),.acc(r108_47),.res(r108_48),.clk(clk),.wout(w108_48));
	PE pe108_49(.x(x49),.w(w108_48),.acc(r108_48),.res(r108_49),.clk(clk),.wout(w108_49));
	PE pe108_50(.x(x50),.w(w108_49),.acc(r108_49),.res(r108_50),.clk(clk),.wout(w108_50));
	PE pe108_51(.x(x51),.w(w108_50),.acc(r108_50),.res(r108_51),.clk(clk),.wout(w108_51));
	PE pe108_52(.x(x52),.w(w108_51),.acc(r108_51),.res(r108_52),.clk(clk),.wout(w108_52));
	PE pe108_53(.x(x53),.w(w108_52),.acc(r108_52),.res(r108_53),.clk(clk),.wout(w108_53));
	PE pe108_54(.x(x54),.w(w108_53),.acc(r108_53),.res(r108_54),.clk(clk),.wout(w108_54));
	PE pe108_55(.x(x55),.w(w108_54),.acc(r108_54),.res(r108_55),.clk(clk),.wout(w108_55));
	PE pe108_56(.x(x56),.w(w108_55),.acc(r108_55),.res(r108_56),.clk(clk),.wout(w108_56));
	PE pe108_57(.x(x57),.w(w108_56),.acc(r108_56),.res(r108_57),.clk(clk),.wout(w108_57));
	PE pe108_58(.x(x58),.w(w108_57),.acc(r108_57),.res(r108_58),.clk(clk),.wout(w108_58));
	PE pe108_59(.x(x59),.w(w108_58),.acc(r108_58),.res(r108_59),.clk(clk),.wout(w108_59));
	PE pe108_60(.x(x60),.w(w108_59),.acc(r108_59),.res(r108_60),.clk(clk),.wout(w108_60));
	PE pe108_61(.x(x61),.w(w108_60),.acc(r108_60),.res(r108_61),.clk(clk),.wout(w108_61));
	PE pe108_62(.x(x62),.w(w108_61),.acc(r108_61),.res(r108_62),.clk(clk),.wout(w108_62));
	PE pe108_63(.x(x63),.w(w108_62),.acc(r108_62),.res(r108_63),.clk(clk),.wout(w108_63));
	PE pe108_64(.x(x64),.w(w108_63),.acc(r108_63),.res(r108_64),.clk(clk),.wout(w108_64));
	PE pe108_65(.x(x65),.w(w108_64),.acc(r108_64),.res(r108_65),.clk(clk),.wout(w108_65));
	PE pe108_66(.x(x66),.w(w108_65),.acc(r108_65),.res(r108_66),.clk(clk),.wout(w108_66));
	PE pe108_67(.x(x67),.w(w108_66),.acc(r108_66),.res(r108_67),.clk(clk),.wout(w108_67));
	PE pe108_68(.x(x68),.w(w108_67),.acc(r108_67),.res(r108_68),.clk(clk),.wout(w108_68));
	PE pe108_69(.x(x69),.w(w108_68),.acc(r108_68),.res(r108_69),.clk(clk),.wout(w108_69));
	PE pe108_70(.x(x70),.w(w108_69),.acc(r108_69),.res(r108_70),.clk(clk),.wout(w108_70));
	PE pe108_71(.x(x71),.w(w108_70),.acc(r108_70),.res(r108_71),.clk(clk),.wout(w108_71));
	PE pe108_72(.x(x72),.w(w108_71),.acc(r108_71),.res(r108_72),.clk(clk),.wout(w108_72));
	PE pe108_73(.x(x73),.w(w108_72),.acc(r108_72),.res(r108_73),.clk(clk),.wout(w108_73));
	PE pe108_74(.x(x74),.w(w108_73),.acc(r108_73),.res(r108_74),.clk(clk),.wout(w108_74));
	PE pe108_75(.x(x75),.w(w108_74),.acc(r108_74),.res(r108_75),.clk(clk),.wout(w108_75));
	PE pe108_76(.x(x76),.w(w108_75),.acc(r108_75),.res(r108_76),.clk(clk),.wout(w108_76));
	PE pe108_77(.x(x77),.w(w108_76),.acc(r108_76),.res(r108_77),.clk(clk),.wout(w108_77));
	PE pe108_78(.x(x78),.w(w108_77),.acc(r108_77),.res(r108_78),.clk(clk),.wout(w108_78));
	PE pe108_79(.x(x79),.w(w108_78),.acc(r108_78),.res(r108_79),.clk(clk),.wout(w108_79));
	PE pe108_80(.x(x80),.w(w108_79),.acc(r108_79),.res(r108_80),.clk(clk),.wout(w108_80));
	PE pe108_81(.x(x81),.w(w108_80),.acc(r108_80),.res(r108_81),.clk(clk),.wout(w108_81));
	PE pe108_82(.x(x82),.w(w108_81),.acc(r108_81),.res(r108_82),.clk(clk),.wout(w108_82));
	PE pe108_83(.x(x83),.w(w108_82),.acc(r108_82),.res(r108_83),.clk(clk),.wout(w108_83));
	PE pe108_84(.x(x84),.w(w108_83),.acc(r108_83),.res(r108_84),.clk(clk),.wout(w108_84));
	PE pe108_85(.x(x85),.w(w108_84),.acc(r108_84),.res(r108_85),.clk(clk),.wout(w108_85));
	PE pe108_86(.x(x86),.w(w108_85),.acc(r108_85),.res(r108_86),.clk(clk),.wout(w108_86));
	PE pe108_87(.x(x87),.w(w108_86),.acc(r108_86),.res(r108_87),.clk(clk),.wout(w108_87));
	PE pe108_88(.x(x88),.w(w108_87),.acc(r108_87),.res(r108_88),.clk(clk),.wout(w108_88));
	PE pe108_89(.x(x89),.w(w108_88),.acc(r108_88),.res(r108_89),.clk(clk),.wout(w108_89));
	PE pe108_90(.x(x90),.w(w108_89),.acc(r108_89),.res(r108_90),.clk(clk),.wout(w108_90));
	PE pe108_91(.x(x91),.w(w108_90),.acc(r108_90),.res(r108_91),.clk(clk),.wout(w108_91));
	PE pe108_92(.x(x92),.w(w108_91),.acc(r108_91),.res(r108_92),.clk(clk),.wout(w108_92));
	PE pe108_93(.x(x93),.w(w108_92),.acc(r108_92),.res(r108_93),.clk(clk),.wout(w108_93));
	PE pe108_94(.x(x94),.w(w108_93),.acc(r108_93),.res(r108_94),.clk(clk),.wout(w108_94));
	PE pe108_95(.x(x95),.w(w108_94),.acc(r108_94),.res(r108_95),.clk(clk),.wout(w108_95));
	PE pe108_96(.x(x96),.w(w108_95),.acc(r108_95),.res(r108_96),.clk(clk),.wout(w108_96));
	PE pe108_97(.x(x97),.w(w108_96),.acc(r108_96),.res(r108_97),.clk(clk),.wout(w108_97));
	PE pe108_98(.x(x98),.w(w108_97),.acc(r108_97),.res(r108_98),.clk(clk),.wout(w108_98));
	PE pe108_99(.x(x99),.w(w108_98),.acc(r108_98),.res(r108_99),.clk(clk),.wout(w108_99));
	PE pe108_100(.x(x100),.w(w108_99),.acc(r108_99),.res(r108_100),.clk(clk),.wout(w108_100));
	PE pe108_101(.x(x101),.w(w108_100),.acc(r108_100),.res(r108_101),.clk(clk),.wout(w108_101));
	PE pe108_102(.x(x102),.w(w108_101),.acc(r108_101),.res(r108_102),.clk(clk),.wout(w108_102));
	PE pe108_103(.x(x103),.w(w108_102),.acc(r108_102),.res(r108_103),.clk(clk),.wout(w108_103));
	PE pe108_104(.x(x104),.w(w108_103),.acc(r108_103),.res(r108_104),.clk(clk),.wout(w108_104));
	PE pe108_105(.x(x105),.w(w108_104),.acc(r108_104),.res(r108_105),.clk(clk),.wout(w108_105));
	PE pe108_106(.x(x106),.w(w108_105),.acc(r108_105),.res(r108_106),.clk(clk),.wout(w108_106));
	PE pe108_107(.x(x107),.w(w108_106),.acc(r108_106),.res(r108_107),.clk(clk),.wout(w108_107));
	PE pe108_108(.x(x108),.w(w108_107),.acc(r108_107),.res(r108_108),.clk(clk),.wout(w108_108));
	PE pe108_109(.x(x109),.w(w108_108),.acc(r108_108),.res(r108_109),.clk(clk),.wout(w108_109));
	PE pe108_110(.x(x110),.w(w108_109),.acc(r108_109),.res(r108_110),.clk(clk),.wout(w108_110));
	PE pe108_111(.x(x111),.w(w108_110),.acc(r108_110),.res(r108_111),.clk(clk),.wout(w108_111));
	PE pe108_112(.x(x112),.w(w108_111),.acc(r108_111),.res(r108_112),.clk(clk),.wout(w108_112));
	PE pe108_113(.x(x113),.w(w108_112),.acc(r108_112),.res(r108_113),.clk(clk),.wout(w108_113));
	PE pe108_114(.x(x114),.w(w108_113),.acc(r108_113),.res(r108_114),.clk(clk),.wout(w108_114));
	PE pe108_115(.x(x115),.w(w108_114),.acc(r108_114),.res(r108_115),.clk(clk),.wout(w108_115));
	PE pe108_116(.x(x116),.w(w108_115),.acc(r108_115),.res(r108_116),.clk(clk),.wout(w108_116));
	PE pe108_117(.x(x117),.w(w108_116),.acc(r108_116),.res(r108_117),.clk(clk),.wout(w108_117));
	PE pe108_118(.x(x118),.w(w108_117),.acc(r108_117),.res(r108_118),.clk(clk),.wout(w108_118));
	PE pe108_119(.x(x119),.w(w108_118),.acc(r108_118),.res(r108_119),.clk(clk),.wout(w108_119));
	PE pe108_120(.x(x120),.w(w108_119),.acc(r108_119),.res(r108_120),.clk(clk),.wout(w108_120));
	PE pe108_121(.x(x121),.w(w108_120),.acc(r108_120),.res(r108_121),.clk(clk),.wout(w108_121));
	PE pe108_122(.x(x122),.w(w108_121),.acc(r108_121),.res(r108_122),.clk(clk),.wout(w108_122));
	PE pe108_123(.x(x123),.w(w108_122),.acc(r108_122),.res(r108_123),.clk(clk),.wout(w108_123));
	PE pe108_124(.x(x124),.w(w108_123),.acc(r108_123),.res(r108_124),.clk(clk),.wout(w108_124));
	PE pe108_125(.x(x125),.w(w108_124),.acc(r108_124),.res(r108_125),.clk(clk),.wout(w108_125));
	PE pe108_126(.x(x126),.w(w108_125),.acc(r108_125),.res(r108_126),.clk(clk),.wout(w108_126));
	PE pe108_127(.x(x127),.w(w108_126),.acc(r108_126),.res(result108),.clk(clk),.wout(weight108));

	PE pe109_0(.x(x0),.w(w109),.acc(32'h0),.res(r109_0),.clk(clk),.wout(w109_0));
	PE pe109_1(.x(x1),.w(w109_0),.acc(r109_0),.res(r109_1),.clk(clk),.wout(w109_1));
	PE pe109_2(.x(x2),.w(w109_1),.acc(r109_1),.res(r109_2),.clk(clk),.wout(w109_2));
	PE pe109_3(.x(x3),.w(w109_2),.acc(r109_2),.res(r109_3),.clk(clk),.wout(w109_3));
	PE pe109_4(.x(x4),.w(w109_3),.acc(r109_3),.res(r109_4),.clk(clk),.wout(w109_4));
	PE pe109_5(.x(x5),.w(w109_4),.acc(r109_4),.res(r109_5),.clk(clk),.wout(w109_5));
	PE pe109_6(.x(x6),.w(w109_5),.acc(r109_5),.res(r109_6),.clk(clk),.wout(w109_6));
	PE pe109_7(.x(x7),.w(w109_6),.acc(r109_6),.res(r109_7),.clk(clk),.wout(w109_7));
	PE pe109_8(.x(x8),.w(w109_7),.acc(r109_7),.res(r109_8),.clk(clk),.wout(w109_8));
	PE pe109_9(.x(x9),.w(w109_8),.acc(r109_8),.res(r109_9),.clk(clk),.wout(w109_9));
	PE pe109_10(.x(x10),.w(w109_9),.acc(r109_9),.res(r109_10),.clk(clk),.wout(w109_10));
	PE pe109_11(.x(x11),.w(w109_10),.acc(r109_10),.res(r109_11),.clk(clk),.wout(w109_11));
	PE pe109_12(.x(x12),.w(w109_11),.acc(r109_11),.res(r109_12),.clk(clk),.wout(w109_12));
	PE pe109_13(.x(x13),.w(w109_12),.acc(r109_12),.res(r109_13),.clk(clk),.wout(w109_13));
	PE pe109_14(.x(x14),.w(w109_13),.acc(r109_13),.res(r109_14),.clk(clk),.wout(w109_14));
	PE pe109_15(.x(x15),.w(w109_14),.acc(r109_14),.res(r109_15),.clk(clk),.wout(w109_15));
	PE pe109_16(.x(x16),.w(w109_15),.acc(r109_15),.res(r109_16),.clk(clk),.wout(w109_16));
	PE pe109_17(.x(x17),.w(w109_16),.acc(r109_16),.res(r109_17),.clk(clk),.wout(w109_17));
	PE pe109_18(.x(x18),.w(w109_17),.acc(r109_17),.res(r109_18),.clk(clk),.wout(w109_18));
	PE pe109_19(.x(x19),.w(w109_18),.acc(r109_18),.res(r109_19),.clk(clk),.wout(w109_19));
	PE pe109_20(.x(x20),.w(w109_19),.acc(r109_19),.res(r109_20),.clk(clk),.wout(w109_20));
	PE pe109_21(.x(x21),.w(w109_20),.acc(r109_20),.res(r109_21),.clk(clk),.wout(w109_21));
	PE pe109_22(.x(x22),.w(w109_21),.acc(r109_21),.res(r109_22),.clk(clk),.wout(w109_22));
	PE pe109_23(.x(x23),.w(w109_22),.acc(r109_22),.res(r109_23),.clk(clk),.wout(w109_23));
	PE pe109_24(.x(x24),.w(w109_23),.acc(r109_23),.res(r109_24),.clk(clk),.wout(w109_24));
	PE pe109_25(.x(x25),.w(w109_24),.acc(r109_24),.res(r109_25),.clk(clk),.wout(w109_25));
	PE pe109_26(.x(x26),.w(w109_25),.acc(r109_25),.res(r109_26),.clk(clk),.wout(w109_26));
	PE pe109_27(.x(x27),.w(w109_26),.acc(r109_26),.res(r109_27),.clk(clk),.wout(w109_27));
	PE pe109_28(.x(x28),.w(w109_27),.acc(r109_27),.res(r109_28),.clk(clk),.wout(w109_28));
	PE pe109_29(.x(x29),.w(w109_28),.acc(r109_28),.res(r109_29),.clk(clk),.wout(w109_29));
	PE pe109_30(.x(x30),.w(w109_29),.acc(r109_29),.res(r109_30),.clk(clk),.wout(w109_30));
	PE pe109_31(.x(x31),.w(w109_30),.acc(r109_30),.res(r109_31),.clk(clk),.wout(w109_31));
	PE pe109_32(.x(x32),.w(w109_31),.acc(r109_31),.res(r109_32),.clk(clk),.wout(w109_32));
	PE pe109_33(.x(x33),.w(w109_32),.acc(r109_32),.res(r109_33),.clk(clk),.wout(w109_33));
	PE pe109_34(.x(x34),.w(w109_33),.acc(r109_33),.res(r109_34),.clk(clk),.wout(w109_34));
	PE pe109_35(.x(x35),.w(w109_34),.acc(r109_34),.res(r109_35),.clk(clk),.wout(w109_35));
	PE pe109_36(.x(x36),.w(w109_35),.acc(r109_35),.res(r109_36),.clk(clk),.wout(w109_36));
	PE pe109_37(.x(x37),.w(w109_36),.acc(r109_36),.res(r109_37),.clk(clk),.wout(w109_37));
	PE pe109_38(.x(x38),.w(w109_37),.acc(r109_37),.res(r109_38),.clk(clk),.wout(w109_38));
	PE pe109_39(.x(x39),.w(w109_38),.acc(r109_38),.res(r109_39),.clk(clk),.wout(w109_39));
	PE pe109_40(.x(x40),.w(w109_39),.acc(r109_39),.res(r109_40),.clk(clk),.wout(w109_40));
	PE pe109_41(.x(x41),.w(w109_40),.acc(r109_40),.res(r109_41),.clk(clk),.wout(w109_41));
	PE pe109_42(.x(x42),.w(w109_41),.acc(r109_41),.res(r109_42),.clk(clk),.wout(w109_42));
	PE pe109_43(.x(x43),.w(w109_42),.acc(r109_42),.res(r109_43),.clk(clk),.wout(w109_43));
	PE pe109_44(.x(x44),.w(w109_43),.acc(r109_43),.res(r109_44),.clk(clk),.wout(w109_44));
	PE pe109_45(.x(x45),.w(w109_44),.acc(r109_44),.res(r109_45),.clk(clk),.wout(w109_45));
	PE pe109_46(.x(x46),.w(w109_45),.acc(r109_45),.res(r109_46),.clk(clk),.wout(w109_46));
	PE pe109_47(.x(x47),.w(w109_46),.acc(r109_46),.res(r109_47),.clk(clk),.wout(w109_47));
	PE pe109_48(.x(x48),.w(w109_47),.acc(r109_47),.res(r109_48),.clk(clk),.wout(w109_48));
	PE pe109_49(.x(x49),.w(w109_48),.acc(r109_48),.res(r109_49),.clk(clk),.wout(w109_49));
	PE pe109_50(.x(x50),.w(w109_49),.acc(r109_49),.res(r109_50),.clk(clk),.wout(w109_50));
	PE pe109_51(.x(x51),.w(w109_50),.acc(r109_50),.res(r109_51),.clk(clk),.wout(w109_51));
	PE pe109_52(.x(x52),.w(w109_51),.acc(r109_51),.res(r109_52),.clk(clk),.wout(w109_52));
	PE pe109_53(.x(x53),.w(w109_52),.acc(r109_52),.res(r109_53),.clk(clk),.wout(w109_53));
	PE pe109_54(.x(x54),.w(w109_53),.acc(r109_53),.res(r109_54),.clk(clk),.wout(w109_54));
	PE pe109_55(.x(x55),.w(w109_54),.acc(r109_54),.res(r109_55),.clk(clk),.wout(w109_55));
	PE pe109_56(.x(x56),.w(w109_55),.acc(r109_55),.res(r109_56),.clk(clk),.wout(w109_56));
	PE pe109_57(.x(x57),.w(w109_56),.acc(r109_56),.res(r109_57),.clk(clk),.wout(w109_57));
	PE pe109_58(.x(x58),.w(w109_57),.acc(r109_57),.res(r109_58),.clk(clk),.wout(w109_58));
	PE pe109_59(.x(x59),.w(w109_58),.acc(r109_58),.res(r109_59),.clk(clk),.wout(w109_59));
	PE pe109_60(.x(x60),.w(w109_59),.acc(r109_59),.res(r109_60),.clk(clk),.wout(w109_60));
	PE pe109_61(.x(x61),.w(w109_60),.acc(r109_60),.res(r109_61),.clk(clk),.wout(w109_61));
	PE pe109_62(.x(x62),.w(w109_61),.acc(r109_61),.res(r109_62),.clk(clk),.wout(w109_62));
	PE pe109_63(.x(x63),.w(w109_62),.acc(r109_62),.res(r109_63),.clk(clk),.wout(w109_63));
	PE pe109_64(.x(x64),.w(w109_63),.acc(r109_63),.res(r109_64),.clk(clk),.wout(w109_64));
	PE pe109_65(.x(x65),.w(w109_64),.acc(r109_64),.res(r109_65),.clk(clk),.wout(w109_65));
	PE pe109_66(.x(x66),.w(w109_65),.acc(r109_65),.res(r109_66),.clk(clk),.wout(w109_66));
	PE pe109_67(.x(x67),.w(w109_66),.acc(r109_66),.res(r109_67),.clk(clk),.wout(w109_67));
	PE pe109_68(.x(x68),.w(w109_67),.acc(r109_67),.res(r109_68),.clk(clk),.wout(w109_68));
	PE pe109_69(.x(x69),.w(w109_68),.acc(r109_68),.res(r109_69),.clk(clk),.wout(w109_69));
	PE pe109_70(.x(x70),.w(w109_69),.acc(r109_69),.res(r109_70),.clk(clk),.wout(w109_70));
	PE pe109_71(.x(x71),.w(w109_70),.acc(r109_70),.res(r109_71),.clk(clk),.wout(w109_71));
	PE pe109_72(.x(x72),.w(w109_71),.acc(r109_71),.res(r109_72),.clk(clk),.wout(w109_72));
	PE pe109_73(.x(x73),.w(w109_72),.acc(r109_72),.res(r109_73),.clk(clk),.wout(w109_73));
	PE pe109_74(.x(x74),.w(w109_73),.acc(r109_73),.res(r109_74),.clk(clk),.wout(w109_74));
	PE pe109_75(.x(x75),.w(w109_74),.acc(r109_74),.res(r109_75),.clk(clk),.wout(w109_75));
	PE pe109_76(.x(x76),.w(w109_75),.acc(r109_75),.res(r109_76),.clk(clk),.wout(w109_76));
	PE pe109_77(.x(x77),.w(w109_76),.acc(r109_76),.res(r109_77),.clk(clk),.wout(w109_77));
	PE pe109_78(.x(x78),.w(w109_77),.acc(r109_77),.res(r109_78),.clk(clk),.wout(w109_78));
	PE pe109_79(.x(x79),.w(w109_78),.acc(r109_78),.res(r109_79),.clk(clk),.wout(w109_79));
	PE pe109_80(.x(x80),.w(w109_79),.acc(r109_79),.res(r109_80),.clk(clk),.wout(w109_80));
	PE pe109_81(.x(x81),.w(w109_80),.acc(r109_80),.res(r109_81),.clk(clk),.wout(w109_81));
	PE pe109_82(.x(x82),.w(w109_81),.acc(r109_81),.res(r109_82),.clk(clk),.wout(w109_82));
	PE pe109_83(.x(x83),.w(w109_82),.acc(r109_82),.res(r109_83),.clk(clk),.wout(w109_83));
	PE pe109_84(.x(x84),.w(w109_83),.acc(r109_83),.res(r109_84),.clk(clk),.wout(w109_84));
	PE pe109_85(.x(x85),.w(w109_84),.acc(r109_84),.res(r109_85),.clk(clk),.wout(w109_85));
	PE pe109_86(.x(x86),.w(w109_85),.acc(r109_85),.res(r109_86),.clk(clk),.wout(w109_86));
	PE pe109_87(.x(x87),.w(w109_86),.acc(r109_86),.res(r109_87),.clk(clk),.wout(w109_87));
	PE pe109_88(.x(x88),.w(w109_87),.acc(r109_87),.res(r109_88),.clk(clk),.wout(w109_88));
	PE pe109_89(.x(x89),.w(w109_88),.acc(r109_88),.res(r109_89),.clk(clk),.wout(w109_89));
	PE pe109_90(.x(x90),.w(w109_89),.acc(r109_89),.res(r109_90),.clk(clk),.wout(w109_90));
	PE pe109_91(.x(x91),.w(w109_90),.acc(r109_90),.res(r109_91),.clk(clk),.wout(w109_91));
	PE pe109_92(.x(x92),.w(w109_91),.acc(r109_91),.res(r109_92),.clk(clk),.wout(w109_92));
	PE pe109_93(.x(x93),.w(w109_92),.acc(r109_92),.res(r109_93),.clk(clk),.wout(w109_93));
	PE pe109_94(.x(x94),.w(w109_93),.acc(r109_93),.res(r109_94),.clk(clk),.wout(w109_94));
	PE pe109_95(.x(x95),.w(w109_94),.acc(r109_94),.res(r109_95),.clk(clk),.wout(w109_95));
	PE pe109_96(.x(x96),.w(w109_95),.acc(r109_95),.res(r109_96),.clk(clk),.wout(w109_96));
	PE pe109_97(.x(x97),.w(w109_96),.acc(r109_96),.res(r109_97),.clk(clk),.wout(w109_97));
	PE pe109_98(.x(x98),.w(w109_97),.acc(r109_97),.res(r109_98),.clk(clk),.wout(w109_98));
	PE pe109_99(.x(x99),.w(w109_98),.acc(r109_98),.res(r109_99),.clk(clk),.wout(w109_99));
	PE pe109_100(.x(x100),.w(w109_99),.acc(r109_99),.res(r109_100),.clk(clk),.wout(w109_100));
	PE pe109_101(.x(x101),.w(w109_100),.acc(r109_100),.res(r109_101),.clk(clk),.wout(w109_101));
	PE pe109_102(.x(x102),.w(w109_101),.acc(r109_101),.res(r109_102),.clk(clk),.wout(w109_102));
	PE pe109_103(.x(x103),.w(w109_102),.acc(r109_102),.res(r109_103),.clk(clk),.wout(w109_103));
	PE pe109_104(.x(x104),.w(w109_103),.acc(r109_103),.res(r109_104),.clk(clk),.wout(w109_104));
	PE pe109_105(.x(x105),.w(w109_104),.acc(r109_104),.res(r109_105),.clk(clk),.wout(w109_105));
	PE pe109_106(.x(x106),.w(w109_105),.acc(r109_105),.res(r109_106),.clk(clk),.wout(w109_106));
	PE pe109_107(.x(x107),.w(w109_106),.acc(r109_106),.res(r109_107),.clk(clk),.wout(w109_107));
	PE pe109_108(.x(x108),.w(w109_107),.acc(r109_107),.res(r109_108),.clk(clk),.wout(w109_108));
	PE pe109_109(.x(x109),.w(w109_108),.acc(r109_108),.res(r109_109),.clk(clk),.wout(w109_109));
	PE pe109_110(.x(x110),.w(w109_109),.acc(r109_109),.res(r109_110),.clk(clk),.wout(w109_110));
	PE pe109_111(.x(x111),.w(w109_110),.acc(r109_110),.res(r109_111),.clk(clk),.wout(w109_111));
	PE pe109_112(.x(x112),.w(w109_111),.acc(r109_111),.res(r109_112),.clk(clk),.wout(w109_112));
	PE pe109_113(.x(x113),.w(w109_112),.acc(r109_112),.res(r109_113),.clk(clk),.wout(w109_113));
	PE pe109_114(.x(x114),.w(w109_113),.acc(r109_113),.res(r109_114),.clk(clk),.wout(w109_114));
	PE pe109_115(.x(x115),.w(w109_114),.acc(r109_114),.res(r109_115),.clk(clk),.wout(w109_115));
	PE pe109_116(.x(x116),.w(w109_115),.acc(r109_115),.res(r109_116),.clk(clk),.wout(w109_116));
	PE pe109_117(.x(x117),.w(w109_116),.acc(r109_116),.res(r109_117),.clk(clk),.wout(w109_117));
	PE pe109_118(.x(x118),.w(w109_117),.acc(r109_117),.res(r109_118),.clk(clk),.wout(w109_118));
	PE pe109_119(.x(x119),.w(w109_118),.acc(r109_118),.res(r109_119),.clk(clk),.wout(w109_119));
	PE pe109_120(.x(x120),.w(w109_119),.acc(r109_119),.res(r109_120),.clk(clk),.wout(w109_120));
	PE pe109_121(.x(x121),.w(w109_120),.acc(r109_120),.res(r109_121),.clk(clk),.wout(w109_121));
	PE pe109_122(.x(x122),.w(w109_121),.acc(r109_121),.res(r109_122),.clk(clk),.wout(w109_122));
	PE pe109_123(.x(x123),.w(w109_122),.acc(r109_122),.res(r109_123),.clk(clk),.wout(w109_123));
	PE pe109_124(.x(x124),.w(w109_123),.acc(r109_123),.res(r109_124),.clk(clk),.wout(w109_124));
	PE pe109_125(.x(x125),.w(w109_124),.acc(r109_124),.res(r109_125),.clk(clk),.wout(w109_125));
	PE pe109_126(.x(x126),.w(w109_125),.acc(r109_125),.res(r109_126),.clk(clk),.wout(w109_126));
	PE pe109_127(.x(x127),.w(w109_126),.acc(r109_126),.res(result109),.clk(clk),.wout(weight109));

	PE pe110_0(.x(x0),.w(w110),.acc(32'h0),.res(r110_0),.clk(clk),.wout(w110_0));
	PE pe110_1(.x(x1),.w(w110_0),.acc(r110_0),.res(r110_1),.clk(clk),.wout(w110_1));
	PE pe110_2(.x(x2),.w(w110_1),.acc(r110_1),.res(r110_2),.clk(clk),.wout(w110_2));
	PE pe110_3(.x(x3),.w(w110_2),.acc(r110_2),.res(r110_3),.clk(clk),.wout(w110_3));
	PE pe110_4(.x(x4),.w(w110_3),.acc(r110_3),.res(r110_4),.clk(clk),.wout(w110_4));
	PE pe110_5(.x(x5),.w(w110_4),.acc(r110_4),.res(r110_5),.clk(clk),.wout(w110_5));
	PE pe110_6(.x(x6),.w(w110_5),.acc(r110_5),.res(r110_6),.clk(clk),.wout(w110_6));
	PE pe110_7(.x(x7),.w(w110_6),.acc(r110_6),.res(r110_7),.clk(clk),.wout(w110_7));
	PE pe110_8(.x(x8),.w(w110_7),.acc(r110_7),.res(r110_8),.clk(clk),.wout(w110_8));
	PE pe110_9(.x(x9),.w(w110_8),.acc(r110_8),.res(r110_9),.clk(clk),.wout(w110_9));
	PE pe110_10(.x(x10),.w(w110_9),.acc(r110_9),.res(r110_10),.clk(clk),.wout(w110_10));
	PE pe110_11(.x(x11),.w(w110_10),.acc(r110_10),.res(r110_11),.clk(clk),.wout(w110_11));
	PE pe110_12(.x(x12),.w(w110_11),.acc(r110_11),.res(r110_12),.clk(clk),.wout(w110_12));
	PE pe110_13(.x(x13),.w(w110_12),.acc(r110_12),.res(r110_13),.clk(clk),.wout(w110_13));
	PE pe110_14(.x(x14),.w(w110_13),.acc(r110_13),.res(r110_14),.clk(clk),.wout(w110_14));
	PE pe110_15(.x(x15),.w(w110_14),.acc(r110_14),.res(r110_15),.clk(clk),.wout(w110_15));
	PE pe110_16(.x(x16),.w(w110_15),.acc(r110_15),.res(r110_16),.clk(clk),.wout(w110_16));
	PE pe110_17(.x(x17),.w(w110_16),.acc(r110_16),.res(r110_17),.clk(clk),.wout(w110_17));
	PE pe110_18(.x(x18),.w(w110_17),.acc(r110_17),.res(r110_18),.clk(clk),.wout(w110_18));
	PE pe110_19(.x(x19),.w(w110_18),.acc(r110_18),.res(r110_19),.clk(clk),.wout(w110_19));
	PE pe110_20(.x(x20),.w(w110_19),.acc(r110_19),.res(r110_20),.clk(clk),.wout(w110_20));
	PE pe110_21(.x(x21),.w(w110_20),.acc(r110_20),.res(r110_21),.clk(clk),.wout(w110_21));
	PE pe110_22(.x(x22),.w(w110_21),.acc(r110_21),.res(r110_22),.clk(clk),.wout(w110_22));
	PE pe110_23(.x(x23),.w(w110_22),.acc(r110_22),.res(r110_23),.clk(clk),.wout(w110_23));
	PE pe110_24(.x(x24),.w(w110_23),.acc(r110_23),.res(r110_24),.clk(clk),.wout(w110_24));
	PE pe110_25(.x(x25),.w(w110_24),.acc(r110_24),.res(r110_25),.clk(clk),.wout(w110_25));
	PE pe110_26(.x(x26),.w(w110_25),.acc(r110_25),.res(r110_26),.clk(clk),.wout(w110_26));
	PE pe110_27(.x(x27),.w(w110_26),.acc(r110_26),.res(r110_27),.clk(clk),.wout(w110_27));
	PE pe110_28(.x(x28),.w(w110_27),.acc(r110_27),.res(r110_28),.clk(clk),.wout(w110_28));
	PE pe110_29(.x(x29),.w(w110_28),.acc(r110_28),.res(r110_29),.clk(clk),.wout(w110_29));
	PE pe110_30(.x(x30),.w(w110_29),.acc(r110_29),.res(r110_30),.clk(clk),.wout(w110_30));
	PE pe110_31(.x(x31),.w(w110_30),.acc(r110_30),.res(r110_31),.clk(clk),.wout(w110_31));
	PE pe110_32(.x(x32),.w(w110_31),.acc(r110_31),.res(r110_32),.clk(clk),.wout(w110_32));
	PE pe110_33(.x(x33),.w(w110_32),.acc(r110_32),.res(r110_33),.clk(clk),.wout(w110_33));
	PE pe110_34(.x(x34),.w(w110_33),.acc(r110_33),.res(r110_34),.clk(clk),.wout(w110_34));
	PE pe110_35(.x(x35),.w(w110_34),.acc(r110_34),.res(r110_35),.clk(clk),.wout(w110_35));
	PE pe110_36(.x(x36),.w(w110_35),.acc(r110_35),.res(r110_36),.clk(clk),.wout(w110_36));
	PE pe110_37(.x(x37),.w(w110_36),.acc(r110_36),.res(r110_37),.clk(clk),.wout(w110_37));
	PE pe110_38(.x(x38),.w(w110_37),.acc(r110_37),.res(r110_38),.clk(clk),.wout(w110_38));
	PE pe110_39(.x(x39),.w(w110_38),.acc(r110_38),.res(r110_39),.clk(clk),.wout(w110_39));
	PE pe110_40(.x(x40),.w(w110_39),.acc(r110_39),.res(r110_40),.clk(clk),.wout(w110_40));
	PE pe110_41(.x(x41),.w(w110_40),.acc(r110_40),.res(r110_41),.clk(clk),.wout(w110_41));
	PE pe110_42(.x(x42),.w(w110_41),.acc(r110_41),.res(r110_42),.clk(clk),.wout(w110_42));
	PE pe110_43(.x(x43),.w(w110_42),.acc(r110_42),.res(r110_43),.clk(clk),.wout(w110_43));
	PE pe110_44(.x(x44),.w(w110_43),.acc(r110_43),.res(r110_44),.clk(clk),.wout(w110_44));
	PE pe110_45(.x(x45),.w(w110_44),.acc(r110_44),.res(r110_45),.clk(clk),.wout(w110_45));
	PE pe110_46(.x(x46),.w(w110_45),.acc(r110_45),.res(r110_46),.clk(clk),.wout(w110_46));
	PE pe110_47(.x(x47),.w(w110_46),.acc(r110_46),.res(r110_47),.clk(clk),.wout(w110_47));
	PE pe110_48(.x(x48),.w(w110_47),.acc(r110_47),.res(r110_48),.clk(clk),.wout(w110_48));
	PE pe110_49(.x(x49),.w(w110_48),.acc(r110_48),.res(r110_49),.clk(clk),.wout(w110_49));
	PE pe110_50(.x(x50),.w(w110_49),.acc(r110_49),.res(r110_50),.clk(clk),.wout(w110_50));
	PE pe110_51(.x(x51),.w(w110_50),.acc(r110_50),.res(r110_51),.clk(clk),.wout(w110_51));
	PE pe110_52(.x(x52),.w(w110_51),.acc(r110_51),.res(r110_52),.clk(clk),.wout(w110_52));
	PE pe110_53(.x(x53),.w(w110_52),.acc(r110_52),.res(r110_53),.clk(clk),.wout(w110_53));
	PE pe110_54(.x(x54),.w(w110_53),.acc(r110_53),.res(r110_54),.clk(clk),.wout(w110_54));
	PE pe110_55(.x(x55),.w(w110_54),.acc(r110_54),.res(r110_55),.clk(clk),.wout(w110_55));
	PE pe110_56(.x(x56),.w(w110_55),.acc(r110_55),.res(r110_56),.clk(clk),.wout(w110_56));
	PE pe110_57(.x(x57),.w(w110_56),.acc(r110_56),.res(r110_57),.clk(clk),.wout(w110_57));
	PE pe110_58(.x(x58),.w(w110_57),.acc(r110_57),.res(r110_58),.clk(clk),.wout(w110_58));
	PE pe110_59(.x(x59),.w(w110_58),.acc(r110_58),.res(r110_59),.clk(clk),.wout(w110_59));
	PE pe110_60(.x(x60),.w(w110_59),.acc(r110_59),.res(r110_60),.clk(clk),.wout(w110_60));
	PE pe110_61(.x(x61),.w(w110_60),.acc(r110_60),.res(r110_61),.clk(clk),.wout(w110_61));
	PE pe110_62(.x(x62),.w(w110_61),.acc(r110_61),.res(r110_62),.clk(clk),.wout(w110_62));
	PE pe110_63(.x(x63),.w(w110_62),.acc(r110_62),.res(r110_63),.clk(clk),.wout(w110_63));
	PE pe110_64(.x(x64),.w(w110_63),.acc(r110_63),.res(r110_64),.clk(clk),.wout(w110_64));
	PE pe110_65(.x(x65),.w(w110_64),.acc(r110_64),.res(r110_65),.clk(clk),.wout(w110_65));
	PE pe110_66(.x(x66),.w(w110_65),.acc(r110_65),.res(r110_66),.clk(clk),.wout(w110_66));
	PE pe110_67(.x(x67),.w(w110_66),.acc(r110_66),.res(r110_67),.clk(clk),.wout(w110_67));
	PE pe110_68(.x(x68),.w(w110_67),.acc(r110_67),.res(r110_68),.clk(clk),.wout(w110_68));
	PE pe110_69(.x(x69),.w(w110_68),.acc(r110_68),.res(r110_69),.clk(clk),.wout(w110_69));
	PE pe110_70(.x(x70),.w(w110_69),.acc(r110_69),.res(r110_70),.clk(clk),.wout(w110_70));
	PE pe110_71(.x(x71),.w(w110_70),.acc(r110_70),.res(r110_71),.clk(clk),.wout(w110_71));
	PE pe110_72(.x(x72),.w(w110_71),.acc(r110_71),.res(r110_72),.clk(clk),.wout(w110_72));
	PE pe110_73(.x(x73),.w(w110_72),.acc(r110_72),.res(r110_73),.clk(clk),.wout(w110_73));
	PE pe110_74(.x(x74),.w(w110_73),.acc(r110_73),.res(r110_74),.clk(clk),.wout(w110_74));
	PE pe110_75(.x(x75),.w(w110_74),.acc(r110_74),.res(r110_75),.clk(clk),.wout(w110_75));
	PE pe110_76(.x(x76),.w(w110_75),.acc(r110_75),.res(r110_76),.clk(clk),.wout(w110_76));
	PE pe110_77(.x(x77),.w(w110_76),.acc(r110_76),.res(r110_77),.clk(clk),.wout(w110_77));
	PE pe110_78(.x(x78),.w(w110_77),.acc(r110_77),.res(r110_78),.clk(clk),.wout(w110_78));
	PE pe110_79(.x(x79),.w(w110_78),.acc(r110_78),.res(r110_79),.clk(clk),.wout(w110_79));
	PE pe110_80(.x(x80),.w(w110_79),.acc(r110_79),.res(r110_80),.clk(clk),.wout(w110_80));
	PE pe110_81(.x(x81),.w(w110_80),.acc(r110_80),.res(r110_81),.clk(clk),.wout(w110_81));
	PE pe110_82(.x(x82),.w(w110_81),.acc(r110_81),.res(r110_82),.clk(clk),.wout(w110_82));
	PE pe110_83(.x(x83),.w(w110_82),.acc(r110_82),.res(r110_83),.clk(clk),.wout(w110_83));
	PE pe110_84(.x(x84),.w(w110_83),.acc(r110_83),.res(r110_84),.clk(clk),.wout(w110_84));
	PE pe110_85(.x(x85),.w(w110_84),.acc(r110_84),.res(r110_85),.clk(clk),.wout(w110_85));
	PE pe110_86(.x(x86),.w(w110_85),.acc(r110_85),.res(r110_86),.clk(clk),.wout(w110_86));
	PE pe110_87(.x(x87),.w(w110_86),.acc(r110_86),.res(r110_87),.clk(clk),.wout(w110_87));
	PE pe110_88(.x(x88),.w(w110_87),.acc(r110_87),.res(r110_88),.clk(clk),.wout(w110_88));
	PE pe110_89(.x(x89),.w(w110_88),.acc(r110_88),.res(r110_89),.clk(clk),.wout(w110_89));
	PE pe110_90(.x(x90),.w(w110_89),.acc(r110_89),.res(r110_90),.clk(clk),.wout(w110_90));
	PE pe110_91(.x(x91),.w(w110_90),.acc(r110_90),.res(r110_91),.clk(clk),.wout(w110_91));
	PE pe110_92(.x(x92),.w(w110_91),.acc(r110_91),.res(r110_92),.clk(clk),.wout(w110_92));
	PE pe110_93(.x(x93),.w(w110_92),.acc(r110_92),.res(r110_93),.clk(clk),.wout(w110_93));
	PE pe110_94(.x(x94),.w(w110_93),.acc(r110_93),.res(r110_94),.clk(clk),.wout(w110_94));
	PE pe110_95(.x(x95),.w(w110_94),.acc(r110_94),.res(r110_95),.clk(clk),.wout(w110_95));
	PE pe110_96(.x(x96),.w(w110_95),.acc(r110_95),.res(r110_96),.clk(clk),.wout(w110_96));
	PE pe110_97(.x(x97),.w(w110_96),.acc(r110_96),.res(r110_97),.clk(clk),.wout(w110_97));
	PE pe110_98(.x(x98),.w(w110_97),.acc(r110_97),.res(r110_98),.clk(clk),.wout(w110_98));
	PE pe110_99(.x(x99),.w(w110_98),.acc(r110_98),.res(r110_99),.clk(clk),.wout(w110_99));
	PE pe110_100(.x(x100),.w(w110_99),.acc(r110_99),.res(r110_100),.clk(clk),.wout(w110_100));
	PE pe110_101(.x(x101),.w(w110_100),.acc(r110_100),.res(r110_101),.clk(clk),.wout(w110_101));
	PE pe110_102(.x(x102),.w(w110_101),.acc(r110_101),.res(r110_102),.clk(clk),.wout(w110_102));
	PE pe110_103(.x(x103),.w(w110_102),.acc(r110_102),.res(r110_103),.clk(clk),.wout(w110_103));
	PE pe110_104(.x(x104),.w(w110_103),.acc(r110_103),.res(r110_104),.clk(clk),.wout(w110_104));
	PE pe110_105(.x(x105),.w(w110_104),.acc(r110_104),.res(r110_105),.clk(clk),.wout(w110_105));
	PE pe110_106(.x(x106),.w(w110_105),.acc(r110_105),.res(r110_106),.clk(clk),.wout(w110_106));
	PE pe110_107(.x(x107),.w(w110_106),.acc(r110_106),.res(r110_107),.clk(clk),.wout(w110_107));
	PE pe110_108(.x(x108),.w(w110_107),.acc(r110_107),.res(r110_108),.clk(clk),.wout(w110_108));
	PE pe110_109(.x(x109),.w(w110_108),.acc(r110_108),.res(r110_109),.clk(clk),.wout(w110_109));
	PE pe110_110(.x(x110),.w(w110_109),.acc(r110_109),.res(r110_110),.clk(clk),.wout(w110_110));
	PE pe110_111(.x(x111),.w(w110_110),.acc(r110_110),.res(r110_111),.clk(clk),.wout(w110_111));
	PE pe110_112(.x(x112),.w(w110_111),.acc(r110_111),.res(r110_112),.clk(clk),.wout(w110_112));
	PE pe110_113(.x(x113),.w(w110_112),.acc(r110_112),.res(r110_113),.clk(clk),.wout(w110_113));
	PE pe110_114(.x(x114),.w(w110_113),.acc(r110_113),.res(r110_114),.clk(clk),.wout(w110_114));
	PE pe110_115(.x(x115),.w(w110_114),.acc(r110_114),.res(r110_115),.clk(clk),.wout(w110_115));
	PE pe110_116(.x(x116),.w(w110_115),.acc(r110_115),.res(r110_116),.clk(clk),.wout(w110_116));
	PE pe110_117(.x(x117),.w(w110_116),.acc(r110_116),.res(r110_117),.clk(clk),.wout(w110_117));
	PE pe110_118(.x(x118),.w(w110_117),.acc(r110_117),.res(r110_118),.clk(clk),.wout(w110_118));
	PE pe110_119(.x(x119),.w(w110_118),.acc(r110_118),.res(r110_119),.clk(clk),.wout(w110_119));
	PE pe110_120(.x(x120),.w(w110_119),.acc(r110_119),.res(r110_120),.clk(clk),.wout(w110_120));
	PE pe110_121(.x(x121),.w(w110_120),.acc(r110_120),.res(r110_121),.clk(clk),.wout(w110_121));
	PE pe110_122(.x(x122),.w(w110_121),.acc(r110_121),.res(r110_122),.clk(clk),.wout(w110_122));
	PE pe110_123(.x(x123),.w(w110_122),.acc(r110_122),.res(r110_123),.clk(clk),.wout(w110_123));
	PE pe110_124(.x(x124),.w(w110_123),.acc(r110_123),.res(r110_124),.clk(clk),.wout(w110_124));
	PE pe110_125(.x(x125),.w(w110_124),.acc(r110_124),.res(r110_125),.clk(clk),.wout(w110_125));
	PE pe110_126(.x(x126),.w(w110_125),.acc(r110_125),.res(r110_126),.clk(clk),.wout(w110_126));
	PE pe110_127(.x(x127),.w(w110_126),.acc(r110_126),.res(result110),.clk(clk),.wout(weight110));

	PE pe111_0(.x(x0),.w(w111),.acc(32'h0),.res(r111_0),.clk(clk),.wout(w111_0));
	PE pe111_1(.x(x1),.w(w111_0),.acc(r111_0),.res(r111_1),.clk(clk),.wout(w111_1));
	PE pe111_2(.x(x2),.w(w111_1),.acc(r111_1),.res(r111_2),.clk(clk),.wout(w111_2));
	PE pe111_3(.x(x3),.w(w111_2),.acc(r111_2),.res(r111_3),.clk(clk),.wout(w111_3));
	PE pe111_4(.x(x4),.w(w111_3),.acc(r111_3),.res(r111_4),.clk(clk),.wout(w111_4));
	PE pe111_5(.x(x5),.w(w111_4),.acc(r111_4),.res(r111_5),.clk(clk),.wout(w111_5));
	PE pe111_6(.x(x6),.w(w111_5),.acc(r111_5),.res(r111_6),.clk(clk),.wout(w111_6));
	PE pe111_7(.x(x7),.w(w111_6),.acc(r111_6),.res(r111_7),.clk(clk),.wout(w111_7));
	PE pe111_8(.x(x8),.w(w111_7),.acc(r111_7),.res(r111_8),.clk(clk),.wout(w111_8));
	PE pe111_9(.x(x9),.w(w111_8),.acc(r111_8),.res(r111_9),.clk(clk),.wout(w111_9));
	PE pe111_10(.x(x10),.w(w111_9),.acc(r111_9),.res(r111_10),.clk(clk),.wout(w111_10));
	PE pe111_11(.x(x11),.w(w111_10),.acc(r111_10),.res(r111_11),.clk(clk),.wout(w111_11));
	PE pe111_12(.x(x12),.w(w111_11),.acc(r111_11),.res(r111_12),.clk(clk),.wout(w111_12));
	PE pe111_13(.x(x13),.w(w111_12),.acc(r111_12),.res(r111_13),.clk(clk),.wout(w111_13));
	PE pe111_14(.x(x14),.w(w111_13),.acc(r111_13),.res(r111_14),.clk(clk),.wout(w111_14));
	PE pe111_15(.x(x15),.w(w111_14),.acc(r111_14),.res(r111_15),.clk(clk),.wout(w111_15));
	PE pe111_16(.x(x16),.w(w111_15),.acc(r111_15),.res(r111_16),.clk(clk),.wout(w111_16));
	PE pe111_17(.x(x17),.w(w111_16),.acc(r111_16),.res(r111_17),.clk(clk),.wout(w111_17));
	PE pe111_18(.x(x18),.w(w111_17),.acc(r111_17),.res(r111_18),.clk(clk),.wout(w111_18));
	PE pe111_19(.x(x19),.w(w111_18),.acc(r111_18),.res(r111_19),.clk(clk),.wout(w111_19));
	PE pe111_20(.x(x20),.w(w111_19),.acc(r111_19),.res(r111_20),.clk(clk),.wout(w111_20));
	PE pe111_21(.x(x21),.w(w111_20),.acc(r111_20),.res(r111_21),.clk(clk),.wout(w111_21));
	PE pe111_22(.x(x22),.w(w111_21),.acc(r111_21),.res(r111_22),.clk(clk),.wout(w111_22));
	PE pe111_23(.x(x23),.w(w111_22),.acc(r111_22),.res(r111_23),.clk(clk),.wout(w111_23));
	PE pe111_24(.x(x24),.w(w111_23),.acc(r111_23),.res(r111_24),.clk(clk),.wout(w111_24));
	PE pe111_25(.x(x25),.w(w111_24),.acc(r111_24),.res(r111_25),.clk(clk),.wout(w111_25));
	PE pe111_26(.x(x26),.w(w111_25),.acc(r111_25),.res(r111_26),.clk(clk),.wout(w111_26));
	PE pe111_27(.x(x27),.w(w111_26),.acc(r111_26),.res(r111_27),.clk(clk),.wout(w111_27));
	PE pe111_28(.x(x28),.w(w111_27),.acc(r111_27),.res(r111_28),.clk(clk),.wout(w111_28));
	PE pe111_29(.x(x29),.w(w111_28),.acc(r111_28),.res(r111_29),.clk(clk),.wout(w111_29));
	PE pe111_30(.x(x30),.w(w111_29),.acc(r111_29),.res(r111_30),.clk(clk),.wout(w111_30));
	PE pe111_31(.x(x31),.w(w111_30),.acc(r111_30),.res(r111_31),.clk(clk),.wout(w111_31));
	PE pe111_32(.x(x32),.w(w111_31),.acc(r111_31),.res(r111_32),.clk(clk),.wout(w111_32));
	PE pe111_33(.x(x33),.w(w111_32),.acc(r111_32),.res(r111_33),.clk(clk),.wout(w111_33));
	PE pe111_34(.x(x34),.w(w111_33),.acc(r111_33),.res(r111_34),.clk(clk),.wout(w111_34));
	PE pe111_35(.x(x35),.w(w111_34),.acc(r111_34),.res(r111_35),.clk(clk),.wout(w111_35));
	PE pe111_36(.x(x36),.w(w111_35),.acc(r111_35),.res(r111_36),.clk(clk),.wout(w111_36));
	PE pe111_37(.x(x37),.w(w111_36),.acc(r111_36),.res(r111_37),.clk(clk),.wout(w111_37));
	PE pe111_38(.x(x38),.w(w111_37),.acc(r111_37),.res(r111_38),.clk(clk),.wout(w111_38));
	PE pe111_39(.x(x39),.w(w111_38),.acc(r111_38),.res(r111_39),.clk(clk),.wout(w111_39));
	PE pe111_40(.x(x40),.w(w111_39),.acc(r111_39),.res(r111_40),.clk(clk),.wout(w111_40));
	PE pe111_41(.x(x41),.w(w111_40),.acc(r111_40),.res(r111_41),.clk(clk),.wout(w111_41));
	PE pe111_42(.x(x42),.w(w111_41),.acc(r111_41),.res(r111_42),.clk(clk),.wout(w111_42));
	PE pe111_43(.x(x43),.w(w111_42),.acc(r111_42),.res(r111_43),.clk(clk),.wout(w111_43));
	PE pe111_44(.x(x44),.w(w111_43),.acc(r111_43),.res(r111_44),.clk(clk),.wout(w111_44));
	PE pe111_45(.x(x45),.w(w111_44),.acc(r111_44),.res(r111_45),.clk(clk),.wout(w111_45));
	PE pe111_46(.x(x46),.w(w111_45),.acc(r111_45),.res(r111_46),.clk(clk),.wout(w111_46));
	PE pe111_47(.x(x47),.w(w111_46),.acc(r111_46),.res(r111_47),.clk(clk),.wout(w111_47));
	PE pe111_48(.x(x48),.w(w111_47),.acc(r111_47),.res(r111_48),.clk(clk),.wout(w111_48));
	PE pe111_49(.x(x49),.w(w111_48),.acc(r111_48),.res(r111_49),.clk(clk),.wout(w111_49));
	PE pe111_50(.x(x50),.w(w111_49),.acc(r111_49),.res(r111_50),.clk(clk),.wout(w111_50));
	PE pe111_51(.x(x51),.w(w111_50),.acc(r111_50),.res(r111_51),.clk(clk),.wout(w111_51));
	PE pe111_52(.x(x52),.w(w111_51),.acc(r111_51),.res(r111_52),.clk(clk),.wout(w111_52));
	PE pe111_53(.x(x53),.w(w111_52),.acc(r111_52),.res(r111_53),.clk(clk),.wout(w111_53));
	PE pe111_54(.x(x54),.w(w111_53),.acc(r111_53),.res(r111_54),.clk(clk),.wout(w111_54));
	PE pe111_55(.x(x55),.w(w111_54),.acc(r111_54),.res(r111_55),.clk(clk),.wout(w111_55));
	PE pe111_56(.x(x56),.w(w111_55),.acc(r111_55),.res(r111_56),.clk(clk),.wout(w111_56));
	PE pe111_57(.x(x57),.w(w111_56),.acc(r111_56),.res(r111_57),.clk(clk),.wout(w111_57));
	PE pe111_58(.x(x58),.w(w111_57),.acc(r111_57),.res(r111_58),.clk(clk),.wout(w111_58));
	PE pe111_59(.x(x59),.w(w111_58),.acc(r111_58),.res(r111_59),.clk(clk),.wout(w111_59));
	PE pe111_60(.x(x60),.w(w111_59),.acc(r111_59),.res(r111_60),.clk(clk),.wout(w111_60));
	PE pe111_61(.x(x61),.w(w111_60),.acc(r111_60),.res(r111_61),.clk(clk),.wout(w111_61));
	PE pe111_62(.x(x62),.w(w111_61),.acc(r111_61),.res(r111_62),.clk(clk),.wout(w111_62));
	PE pe111_63(.x(x63),.w(w111_62),.acc(r111_62),.res(r111_63),.clk(clk),.wout(w111_63));
	PE pe111_64(.x(x64),.w(w111_63),.acc(r111_63),.res(r111_64),.clk(clk),.wout(w111_64));
	PE pe111_65(.x(x65),.w(w111_64),.acc(r111_64),.res(r111_65),.clk(clk),.wout(w111_65));
	PE pe111_66(.x(x66),.w(w111_65),.acc(r111_65),.res(r111_66),.clk(clk),.wout(w111_66));
	PE pe111_67(.x(x67),.w(w111_66),.acc(r111_66),.res(r111_67),.clk(clk),.wout(w111_67));
	PE pe111_68(.x(x68),.w(w111_67),.acc(r111_67),.res(r111_68),.clk(clk),.wout(w111_68));
	PE pe111_69(.x(x69),.w(w111_68),.acc(r111_68),.res(r111_69),.clk(clk),.wout(w111_69));
	PE pe111_70(.x(x70),.w(w111_69),.acc(r111_69),.res(r111_70),.clk(clk),.wout(w111_70));
	PE pe111_71(.x(x71),.w(w111_70),.acc(r111_70),.res(r111_71),.clk(clk),.wout(w111_71));
	PE pe111_72(.x(x72),.w(w111_71),.acc(r111_71),.res(r111_72),.clk(clk),.wout(w111_72));
	PE pe111_73(.x(x73),.w(w111_72),.acc(r111_72),.res(r111_73),.clk(clk),.wout(w111_73));
	PE pe111_74(.x(x74),.w(w111_73),.acc(r111_73),.res(r111_74),.clk(clk),.wout(w111_74));
	PE pe111_75(.x(x75),.w(w111_74),.acc(r111_74),.res(r111_75),.clk(clk),.wout(w111_75));
	PE pe111_76(.x(x76),.w(w111_75),.acc(r111_75),.res(r111_76),.clk(clk),.wout(w111_76));
	PE pe111_77(.x(x77),.w(w111_76),.acc(r111_76),.res(r111_77),.clk(clk),.wout(w111_77));
	PE pe111_78(.x(x78),.w(w111_77),.acc(r111_77),.res(r111_78),.clk(clk),.wout(w111_78));
	PE pe111_79(.x(x79),.w(w111_78),.acc(r111_78),.res(r111_79),.clk(clk),.wout(w111_79));
	PE pe111_80(.x(x80),.w(w111_79),.acc(r111_79),.res(r111_80),.clk(clk),.wout(w111_80));
	PE pe111_81(.x(x81),.w(w111_80),.acc(r111_80),.res(r111_81),.clk(clk),.wout(w111_81));
	PE pe111_82(.x(x82),.w(w111_81),.acc(r111_81),.res(r111_82),.clk(clk),.wout(w111_82));
	PE pe111_83(.x(x83),.w(w111_82),.acc(r111_82),.res(r111_83),.clk(clk),.wout(w111_83));
	PE pe111_84(.x(x84),.w(w111_83),.acc(r111_83),.res(r111_84),.clk(clk),.wout(w111_84));
	PE pe111_85(.x(x85),.w(w111_84),.acc(r111_84),.res(r111_85),.clk(clk),.wout(w111_85));
	PE pe111_86(.x(x86),.w(w111_85),.acc(r111_85),.res(r111_86),.clk(clk),.wout(w111_86));
	PE pe111_87(.x(x87),.w(w111_86),.acc(r111_86),.res(r111_87),.clk(clk),.wout(w111_87));
	PE pe111_88(.x(x88),.w(w111_87),.acc(r111_87),.res(r111_88),.clk(clk),.wout(w111_88));
	PE pe111_89(.x(x89),.w(w111_88),.acc(r111_88),.res(r111_89),.clk(clk),.wout(w111_89));
	PE pe111_90(.x(x90),.w(w111_89),.acc(r111_89),.res(r111_90),.clk(clk),.wout(w111_90));
	PE pe111_91(.x(x91),.w(w111_90),.acc(r111_90),.res(r111_91),.clk(clk),.wout(w111_91));
	PE pe111_92(.x(x92),.w(w111_91),.acc(r111_91),.res(r111_92),.clk(clk),.wout(w111_92));
	PE pe111_93(.x(x93),.w(w111_92),.acc(r111_92),.res(r111_93),.clk(clk),.wout(w111_93));
	PE pe111_94(.x(x94),.w(w111_93),.acc(r111_93),.res(r111_94),.clk(clk),.wout(w111_94));
	PE pe111_95(.x(x95),.w(w111_94),.acc(r111_94),.res(r111_95),.clk(clk),.wout(w111_95));
	PE pe111_96(.x(x96),.w(w111_95),.acc(r111_95),.res(r111_96),.clk(clk),.wout(w111_96));
	PE pe111_97(.x(x97),.w(w111_96),.acc(r111_96),.res(r111_97),.clk(clk),.wout(w111_97));
	PE pe111_98(.x(x98),.w(w111_97),.acc(r111_97),.res(r111_98),.clk(clk),.wout(w111_98));
	PE pe111_99(.x(x99),.w(w111_98),.acc(r111_98),.res(r111_99),.clk(clk),.wout(w111_99));
	PE pe111_100(.x(x100),.w(w111_99),.acc(r111_99),.res(r111_100),.clk(clk),.wout(w111_100));
	PE pe111_101(.x(x101),.w(w111_100),.acc(r111_100),.res(r111_101),.clk(clk),.wout(w111_101));
	PE pe111_102(.x(x102),.w(w111_101),.acc(r111_101),.res(r111_102),.clk(clk),.wout(w111_102));
	PE pe111_103(.x(x103),.w(w111_102),.acc(r111_102),.res(r111_103),.clk(clk),.wout(w111_103));
	PE pe111_104(.x(x104),.w(w111_103),.acc(r111_103),.res(r111_104),.clk(clk),.wout(w111_104));
	PE pe111_105(.x(x105),.w(w111_104),.acc(r111_104),.res(r111_105),.clk(clk),.wout(w111_105));
	PE pe111_106(.x(x106),.w(w111_105),.acc(r111_105),.res(r111_106),.clk(clk),.wout(w111_106));
	PE pe111_107(.x(x107),.w(w111_106),.acc(r111_106),.res(r111_107),.clk(clk),.wout(w111_107));
	PE pe111_108(.x(x108),.w(w111_107),.acc(r111_107),.res(r111_108),.clk(clk),.wout(w111_108));
	PE pe111_109(.x(x109),.w(w111_108),.acc(r111_108),.res(r111_109),.clk(clk),.wout(w111_109));
	PE pe111_110(.x(x110),.w(w111_109),.acc(r111_109),.res(r111_110),.clk(clk),.wout(w111_110));
	PE pe111_111(.x(x111),.w(w111_110),.acc(r111_110),.res(r111_111),.clk(clk),.wout(w111_111));
	PE pe111_112(.x(x112),.w(w111_111),.acc(r111_111),.res(r111_112),.clk(clk),.wout(w111_112));
	PE pe111_113(.x(x113),.w(w111_112),.acc(r111_112),.res(r111_113),.clk(clk),.wout(w111_113));
	PE pe111_114(.x(x114),.w(w111_113),.acc(r111_113),.res(r111_114),.clk(clk),.wout(w111_114));
	PE pe111_115(.x(x115),.w(w111_114),.acc(r111_114),.res(r111_115),.clk(clk),.wout(w111_115));
	PE pe111_116(.x(x116),.w(w111_115),.acc(r111_115),.res(r111_116),.clk(clk),.wout(w111_116));
	PE pe111_117(.x(x117),.w(w111_116),.acc(r111_116),.res(r111_117),.clk(clk),.wout(w111_117));
	PE pe111_118(.x(x118),.w(w111_117),.acc(r111_117),.res(r111_118),.clk(clk),.wout(w111_118));
	PE pe111_119(.x(x119),.w(w111_118),.acc(r111_118),.res(r111_119),.clk(clk),.wout(w111_119));
	PE pe111_120(.x(x120),.w(w111_119),.acc(r111_119),.res(r111_120),.clk(clk),.wout(w111_120));
	PE pe111_121(.x(x121),.w(w111_120),.acc(r111_120),.res(r111_121),.clk(clk),.wout(w111_121));
	PE pe111_122(.x(x122),.w(w111_121),.acc(r111_121),.res(r111_122),.clk(clk),.wout(w111_122));
	PE pe111_123(.x(x123),.w(w111_122),.acc(r111_122),.res(r111_123),.clk(clk),.wout(w111_123));
	PE pe111_124(.x(x124),.w(w111_123),.acc(r111_123),.res(r111_124),.clk(clk),.wout(w111_124));
	PE pe111_125(.x(x125),.w(w111_124),.acc(r111_124),.res(r111_125),.clk(clk),.wout(w111_125));
	PE pe111_126(.x(x126),.w(w111_125),.acc(r111_125),.res(r111_126),.clk(clk),.wout(w111_126));
	PE pe111_127(.x(x127),.w(w111_126),.acc(r111_126),.res(result111),.clk(clk),.wout(weight111));

	PE pe112_0(.x(x0),.w(w112),.acc(32'h0),.res(r112_0),.clk(clk),.wout(w112_0));
	PE pe112_1(.x(x1),.w(w112_0),.acc(r112_0),.res(r112_1),.clk(clk),.wout(w112_1));
	PE pe112_2(.x(x2),.w(w112_1),.acc(r112_1),.res(r112_2),.clk(clk),.wout(w112_2));
	PE pe112_3(.x(x3),.w(w112_2),.acc(r112_2),.res(r112_3),.clk(clk),.wout(w112_3));
	PE pe112_4(.x(x4),.w(w112_3),.acc(r112_3),.res(r112_4),.clk(clk),.wout(w112_4));
	PE pe112_5(.x(x5),.w(w112_4),.acc(r112_4),.res(r112_5),.clk(clk),.wout(w112_5));
	PE pe112_6(.x(x6),.w(w112_5),.acc(r112_5),.res(r112_6),.clk(clk),.wout(w112_6));
	PE pe112_7(.x(x7),.w(w112_6),.acc(r112_6),.res(r112_7),.clk(clk),.wout(w112_7));
	PE pe112_8(.x(x8),.w(w112_7),.acc(r112_7),.res(r112_8),.clk(clk),.wout(w112_8));
	PE pe112_9(.x(x9),.w(w112_8),.acc(r112_8),.res(r112_9),.clk(clk),.wout(w112_9));
	PE pe112_10(.x(x10),.w(w112_9),.acc(r112_9),.res(r112_10),.clk(clk),.wout(w112_10));
	PE pe112_11(.x(x11),.w(w112_10),.acc(r112_10),.res(r112_11),.clk(clk),.wout(w112_11));
	PE pe112_12(.x(x12),.w(w112_11),.acc(r112_11),.res(r112_12),.clk(clk),.wout(w112_12));
	PE pe112_13(.x(x13),.w(w112_12),.acc(r112_12),.res(r112_13),.clk(clk),.wout(w112_13));
	PE pe112_14(.x(x14),.w(w112_13),.acc(r112_13),.res(r112_14),.clk(clk),.wout(w112_14));
	PE pe112_15(.x(x15),.w(w112_14),.acc(r112_14),.res(r112_15),.clk(clk),.wout(w112_15));
	PE pe112_16(.x(x16),.w(w112_15),.acc(r112_15),.res(r112_16),.clk(clk),.wout(w112_16));
	PE pe112_17(.x(x17),.w(w112_16),.acc(r112_16),.res(r112_17),.clk(clk),.wout(w112_17));
	PE pe112_18(.x(x18),.w(w112_17),.acc(r112_17),.res(r112_18),.clk(clk),.wout(w112_18));
	PE pe112_19(.x(x19),.w(w112_18),.acc(r112_18),.res(r112_19),.clk(clk),.wout(w112_19));
	PE pe112_20(.x(x20),.w(w112_19),.acc(r112_19),.res(r112_20),.clk(clk),.wout(w112_20));
	PE pe112_21(.x(x21),.w(w112_20),.acc(r112_20),.res(r112_21),.clk(clk),.wout(w112_21));
	PE pe112_22(.x(x22),.w(w112_21),.acc(r112_21),.res(r112_22),.clk(clk),.wout(w112_22));
	PE pe112_23(.x(x23),.w(w112_22),.acc(r112_22),.res(r112_23),.clk(clk),.wout(w112_23));
	PE pe112_24(.x(x24),.w(w112_23),.acc(r112_23),.res(r112_24),.clk(clk),.wout(w112_24));
	PE pe112_25(.x(x25),.w(w112_24),.acc(r112_24),.res(r112_25),.clk(clk),.wout(w112_25));
	PE pe112_26(.x(x26),.w(w112_25),.acc(r112_25),.res(r112_26),.clk(clk),.wout(w112_26));
	PE pe112_27(.x(x27),.w(w112_26),.acc(r112_26),.res(r112_27),.clk(clk),.wout(w112_27));
	PE pe112_28(.x(x28),.w(w112_27),.acc(r112_27),.res(r112_28),.clk(clk),.wout(w112_28));
	PE pe112_29(.x(x29),.w(w112_28),.acc(r112_28),.res(r112_29),.clk(clk),.wout(w112_29));
	PE pe112_30(.x(x30),.w(w112_29),.acc(r112_29),.res(r112_30),.clk(clk),.wout(w112_30));
	PE pe112_31(.x(x31),.w(w112_30),.acc(r112_30),.res(r112_31),.clk(clk),.wout(w112_31));
	PE pe112_32(.x(x32),.w(w112_31),.acc(r112_31),.res(r112_32),.clk(clk),.wout(w112_32));
	PE pe112_33(.x(x33),.w(w112_32),.acc(r112_32),.res(r112_33),.clk(clk),.wout(w112_33));
	PE pe112_34(.x(x34),.w(w112_33),.acc(r112_33),.res(r112_34),.clk(clk),.wout(w112_34));
	PE pe112_35(.x(x35),.w(w112_34),.acc(r112_34),.res(r112_35),.clk(clk),.wout(w112_35));
	PE pe112_36(.x(x36),.w(w112_35),.acc(r112_35),.res(r112_36),.clk(clk),.wout(w112_36));
	PE pe112_37(.x(x37),.w(w112_36),.acc(r112_36),.res(r112_37),.clk(clk),.wout(w112_37));
	PE pe112_38(.x(x38),.w(w112_37),.acc(r112_37),.res(r112_38),.clk(clk),.wout(w112_38));
	PE pe112_39(.x(x39),.w(w112_38),.acc(r112_38),.res(r112_39),.clk(clk),.wout(w112_39));
	PE pe112_40(.x(x40),.w(w112_39),.acc(r112_39),.res(r112_40),.clk(clk),.wout(w112_40));
	PE pe112_41(.x(x41),.w(w112_40),.acc(r112_40),.res(r112_41),.clk(clk),.wout(w112_41));
	PE pe112_42(.x(x42),.w(w112_41),.acc(r112_41),.res(r112_42),.clk(clk),.wout(w112_42));
	PE pe112_43(.x(x43),.w(w112_42),.acc(r112_42),.res(r112_43),.clk(clk),.wout(w112_43));
	PE pe112_44(.x(x44),.w(w112_43),.acc(r112_43),.res(r112_44),.clk(clk),.wout(w112_44));
	PE pe112_45(.x(x45),.w(w112_44),.acc(r112_44),.res(r112_45),.clk(clk),.wout(w112_45));
	PE pe112_46(.x(x46),.w(w112_45),.acc(r112_45),.res(r112_46),.clk(clk),.wout(w112_46));
	PE pe112_47(.x(x47),.w(w112_46),.acc(r112_46),.res(r112_47),.clk(clk),.wout(w112_47));
	PE pe112_48(.x(x48),.w(w112_47),.acc(r112_47),.res(r112_48),.clk(clk),.wout(w112_48));
	PE pe112_49(.x(x49),.w(w112_48),.acc(r112_48),.res(r112_49),.clk(clk),.wout(w112_49));
	PE pe112_50(.x(x50),.w(w112_49),.acc(r112_49),.res(r112_50),.clk(clk),.wout(w112_50));
	PE pe112_51(.x(x51),.w(w112_50),.acc(r112_50),.res(r112_51),.clk(clk),.wout(w112_51));
	PE pe112_52(.x(x52),.w(w112_51),.acc(r112_51),.res(r112_52),.clk(clk),.wout(w112_52));
	PE pe112_53(.x(x53),.w(w112_52),.acc(r112_52),.res(r112_53),.clk(clk),.wout(w112_53));
	PE pe112_54(.x(x54),.w(w112_53),.acc(r112_53),.res(r112_54),.clk(clk),.wout(w112_54));
	PE pe112_55(.x(x55),.w(w112_54),.acc(r112_54),.res(r112_55),.clk(clk),.wout(w112_55));
	PE pe112_56(.x(x56),.w(w112_55),.acc(r112_55),.res(r112_56),.clk(clk),.wout(w112_56));
	PE pe112_57(.x(x57),.w(w112_56),.acc(r112_56),.res(r112_57),.clk(clk),.wout(w112_57));
	PE pe112_58(.x(x58),.w(w112_57),.acc(r112_57),.res(r112_58),.clk(clk),.wout(w112_58));
	PE pe112_59(.x(x59),.w(w112_58),.acc(r112_58),.res(r112_59),.clk(clk),.wout(w112_59));
	PE pe112_60(.x(x60),.w(w112_59),.acc(r112_59),.res(r112_60),.clk(clk),.wout(w112_60));
	PE pe112_61(.x(x61),.w(w112_60),.acc(r112_60),.res(r112_61),.clk(clk),.wout(w112_61));
	PE pe112_62(.x(x62),.w(w112_61),.acc(r112_61),.res(r112_62),.clk(clk),.wout(w112_62));
	PE pe112_63(.x(x63),.w(w112_62),.acc(r112_62),.res(r112_63),.clk(clk),.wout(w112_63));
	PE pe112_64(.x(x64),.w(w112_63),.acc(r112_63),.res(r112_64),.clk(clk),.wout(w112_64));
	PE pe112_65(.x(x65),.w(w112_64),.acc(r112_64),.res(r112_65),.clk(clk),.wout(w112_65));
	PE pe112_66(.x(x66),.w(w112_65),.acc(r112_65),.res(r112_66),.clk(clk),.wout(w112_66));
	PE pe112_67(.x(x67),.w(w112_66),.acc(r112_66),.res(r112_67),.clk(clk),.wout(w112_67));
	PE pe112_68(.x(x68),.w(w112_67),.acc(r112_67),.res(r112_68),.clk(clk),.wout(w112_68));
	PE pe112_69(.x(x69),.w(w112_68),.acc(r112_68),.res(r112_69),.clk(clk),.wout(w112_69));
	PE pe112_70(.x(x70),.w(w112_69),.acc(r112_69),.res(r112_70),.clk(clk),.wout(w112_70));
	PE pe112_71(.x(x71),.w(w112_70),.acc(r112_70),.res(r112_71),.clk(clk),.wout(w112_71));
	PE pe112_72(.x(x72),.w(w112_71),.acc(r112_71),.res(r112_72),.clk(clk),.wout(w112_72));
	PE pe112_73(.x(x73),.w(w112_72),.acc(r112_72),.res(r112_73),.clk(clk),.wout(w112_73));
	PE pe112_74(.x(x74),.w(w112_73),.acc(r112_73),.res(r112_74),.clk(clk),.wout(w112_74));
	PE pe112_75(.x(x75),.w(w112_74),.acc(r112_74),.res(r112_75),.clk(clk),.wout(w112_75));
	PE pe112_76(.x(x76),.w(w112_75),.acc(r112_75),.res(r112_76),.clk(clk),.wout(w112_76));
	PE pe112_77(.x(x77),.w(w112_76),.acc(r112_76),.res(r112_77),.clk(clk),.wout(w112_77));
	PE pe112_78(.x(x78),.w(w112_77),.acc(r112_77),.res(r112_78),.clk(clk),.wout(w112_78));
	PE pe112_79(.x(x79),.w(w112_78),.acc(r112_78),.res(r112_79),.clk(clk),.wout(w112_79));
	PE pe112_80(.x(x80),.w(w112_79),.acc(r112_79),.res(r112_80),.clk(clk),.wout(w112_80));
	PE pe112_81(.x(x81),.w(w112_80),.acc(r112_80),.res(r112_81),.clk(clk),.wout(w112_81));
	PE pe112_82(.x(x82),.w(w112_81),.acc(r112_81),.res(r112_82),.clk(clk),.wout(w112_82));
	PE pe112_83(.x(x83),.w(w112_82),.acc(r112_82),.res(r112_83),.clk(clk),.wout(w112_83));
	PE pe112_84(.x(x84),.w(w112_83),.acc(r112_83),.res(r112_84),.clk(clk),.wout(w112_84));
	PE pe112_85(.x(x85),.w(w112_84),.acc(r112_84),.res(r112_85),.clk(clk),.wout(w112_85));
	PE pe112_86(.x(x86),.w(w112_85),.acc(r112_85),.res(r112_86),.clk(clk),.wout(w112_86));
	PE pe112_87(.x(x87),.w(w112_86),.acc(r112_86),.res(r112_87),.clk(clk),.wout(w112_87));
	PE pe112_88(.x(x88),.w(w112_87),.acc(r112_87),.res(r112_88),.clk(clk),.wout(w112_88));
	PE pe112_89(.x(x89),.w(w112_88),.acc(r112_88),.res(r112_89),.clk(clk),.wout(w112_89));
	PE pe112_90(.x(x90),.w(w112_89),.acc(r112_89),.res(r112_90),.clk(clk),.wout(w112_90));
	PE pe112_91(.x(x91),.w(w112_90),.acc(r112_90),.res(r112_91),.clk(clk),.wout(w112_91));
	PE pe112_92(.x(x92),.w(w112_91),.acc(r112_91),.res(r112_92),.clk(clk),.wout(w112_92));
	PE pe112_93(.x(x93),.w(w112_92),.acc(r112_92),.res(r112_93),.clk(clk),.wout(w112_93));
	PE pe112_94(.x(x94),.w(w112_93),.acc(r112_93),.res(r112_94),.clk(clk),.wout(w112_94));
	PE pe112_95(.x(x95),.w(w112_94),.acc(r112_94),.res(r112_95),.clk(clk),.wout(w112_95));
	PE pe112_96(.x(x96),.w(w112_95),.acc(r112_95),.res(r112_96),.clk(clk),.wout(w112_96));
	PE pe112_97(.x(x97),.w(w112_96),.acc(r112_96),.res(r112_97),.clk(clk),.wout(w112_97));
	PE pe112_98(.x(x98),.w(w112_97),.acc(r112_97),.res(r112_98),.clk(clk),.wout(w112_98));
	PE pe112_99(.x(x99),.w(w112_98),.acc(r112_98),.res(r112_99),.clk(clk),.wout(w112_99));
	PE pe112_100(.x(x100),.w(w112_99),.acc(r112_99),.res(r112_100),.clk(clk),.wout(w112_100));
	PE pe112_101(.x(x101),.w(w112_100),.acc(r112_100),.res(r112_101),.clk(clk),.wout(w112_101));
	PE pe112_102(.x(x102),.w(w112_101),.acc(r112_101),.res(r112_102),.clk(clk),.wout(w112_102));
	PE pe112_103(.x(x103),.w(w112_102),.acc(r112_102),.res(r112_103),.clk(clk),.wout(w112_103));
	PE pe112_104(.x(x104),.w(w112_103),.acc(r112_103),.res(r112_104),.clk(clk),.wout(w112_104));
	PE pe112_105(.x(x105),.w(w112_104),.acc(r112_104),.res(r112_105),.clk(clk),.wout(w112_105));
	PE pe112_106(.x(x106),.w(w112_105),.acc(r112_105),.res(r112_106),.clk(clk),.wout(w112_106));
	PE pe112_107(.x(x107),.w(w112_106),.acc(r112_106),.res(r112_107),.clk(clk),.wout(w112_107));
	PE pe112_108(.x(x108),.w(w112_107),.acc(r112_107),.res(r112_108),.clk(clk),.wout(w112_108));
	PE pe112_109(.x(x109),.w(w112_108),.acc(r112_108),.res(r112_109),.clk(clk),.wout(w112_109));
	PE pe112_110(.x(x110),.w(w112_109),.acc(r112_109),.res(r112_110),.clk(clk),.wout(w112_110));
	PE pe112_111(.x(x111),.w(w112_110),.acc(r112_110),.res(r112_111),.clk(clk),.wout(w112_111));
	PE pe112_112(.x(x112),.w(w112_111),.acc(r112_111),.res(r112_112),.clk(clk),.wout(w112_112));
	PE pe112_113(.x(x113),.w(w112_112),.acc(r112_112),.res(r112_113),.clk(clk),.wout(w112_113));
	PE pe112_114(.x(x114),.w(w112_113),.acc(r112_113),.res(r112_114),.clk(clk),.wout(w112_114));
	PE pe112_115(.x(x115),.w(w112_114),.acc(r112_114),.res(r112_115),.clk(clk),.wout(w112_115));
	PE pe112_116(.x(x116),.w(w112_115),.acc(r112_115),.res(r112_116),.clk(clk),.wout(w112_116));
	PE pe112_117(.x(x117),.w(w112_116),.acc(r112_116),.res(r112_117),.clk(clk),.wout(w112_117));
	PE pe112_118(.x(x118),.w(w112_117),.acc(r112_117),.res(r112_118),.clk(clk),.wout(w112_118));
	PE pe112_119(.x(x119),.w(w112_118),.acc(r112_118),.res(r112_119),.clk(clk),.wout(w112_119));
	PE pe112_120(.x(x120),.w(w112_119),.acc(r112_119),.res(r112_120),.clk(clk),.wout(w112_120));
	PE pe112_121(.x(x121),.w(w112_120),.acc(r112_120),.res(r112_121),.clk(clk),.wout(w112_121));
	PE pe112_122(.x(x122),.w(w112_121),.acc(r112_121),.res(r112_122),.clk(clk),.wout(w112_122));
	PE pe112_123(.x(x123),.w(w112_122),.acc(r112_122),.res(r112_123),.clk(clk),.wout(w112_123));
	PE pe112_124(.x(x124),.w(w112_123),.acc(r112_123),.res(r112_124),.clk(clk),.wout(w112_124));
	PE pe112_125(.x(x125),.w(w112_124),.acc(r112_124),.res(r112_125),.clk(clk),.wout(w112_125));
	PE pe112_126(.x(x126),.w(w112_125),.acc(r112_125),.res(r112_126),.clk(clk),.wout(w112_126));
	PE pe112_127(.x(x127),.w(w112_126),.acc(r112_126),.res(result112),.clk(clk),.wout(weight112));

	PE pe113_0(.x(x0),.w(w113),.acc(32'h0),.res(r113_0),.clk(clk),.wout(w113_0));
	PE pe113_1(.x(x1),.w(w113_0),.acc(r113_0),.res(r113_1),.clk(clk),.wout(w113_1));
	PE pe113_2(.x(x2),.w(w113_1),.acc(r113_1),.res(r113_2),.clk(clk),.wout(w113_2));
	PE pe113_3(.x(x3),.w(w113_2),.acc(r113_2),.res(r113_3),.clk(clk),.wout(w113_3));
	PE pe113_4(.x(x4),.w(w113_3),.acc(r113_3),.res(r113_4),.clk(clk),.wout(w113_4));
	PE pe113_5(.x(x5),.w(w113_4),.acc(r113_4),.res(r113_5),.clk(clk),.wout(w113_5));
	PE pe113_6(.x(x6),.w(w113_5),.acc(r113_5),.res(r113_6),.clk(clk),.wout(w113_6));
	PE pe113_7(.x(x7),.w(w113_6),.acc(r113_6),.res(r113_7),.clk(clk),.wout(w113_7));
	PE pe113_8(.x(x8),.w(w113_7),.acc(r113_7),.res(r113_8),.clk(clk),.wout(w113_8));
	PE pe113_9(.x(x9),.w(w113_8),.acc(r113_8),.res(r113_9),.clk(clk),.wout(w113_9));
	PE pe113_10(.x(x10),.w(w113_9),.acc(r113_9),.res(r113_10),.clk(clk),.wout(w113_10));
	PE pe113_11(.x(x11),.w(w113_10),.acc(r113_10),.res(r113_11),.clk(clk),.wout(w113_11));
	PE pe113_12(.x(x12),.w(w113_11),.acc(r113_11),.res(r113_12),.clk(clk),.wout(w113_12));
	PE pe113_13(.x(x13),.w(w113_12),.acc(r113_12),.res(r113_13),.clk(clk),.wout(w113_13));
	PE pe113_14(.x(x14),.w(w113_13),.acc(r113_13),.res(r113_14),.clk(clk),.wout(w113_14));
	PE pe113_15(.x(x15),.w(w113_14),.acc(r113_14),.res(r113_15),.clk(clk),.wout(w113_15));
	PE pe113_16(.x(x16),.w(w113_15),.acc(r113_15),.res(r113_16),.clk(clk),.wout(w113_16));
	PE pe113_17(.x(x17),.w(w113_16),.acc(r113_16),.res(r113_17),.clk(clk),.wout(w113_17));
	PE pe113_18(.x(x18),.w(w113_17),.acc(r113_17),.res(r113_18),.clk(clk),.wout(w113_18));
	PE pe113_19(.x(x19),.w(w113_18),.acc(r113_18),.res(r113_19),.clk(clk),.wout(w113_19));
	PE pe113_20(.x(x20),.w(w113_19),.acc(r113_19),.res(r113_20),.clk(clk),.wout(w113_20));
	PE pe113_21(.x(x21),.w(w113_20),.acc(r113_20),.res(r113_21),.clk(clk),.wout(w113_21));
	PE pe113_22(.x(x22),.w(w113_21),.acc(r113_21),.res(r113_22),.clk(clk),.wout(w113_22));
	PE pe113_23(.x(x23),.w(w113_22),.acc(r113_22),.res(r113_23),.clk(clk),.wout(w113_23));
	PE pe113_24(.x(x24),.w(w113_23),.acc(r113_23),.res(r113_24),.clk(clk),.wout(w113_24));
	PE pe113_25(.x(x25),.w(w113_24),.acc(r113_24),.res(r113_25),.clk(clk),.wout(w113_25));
	PE pe113_26(.x(x26),.w(w113_25),.acc(r113_25),.res(r113_26),.clk(clk),.wout(w113_26));
	PE pe113_27(.x(x27),.w(w113_26),.acc(r113_26),.res(r113_27),.clk(clk),.wout(w113_27));
	PE pe113_28(.x(x28),.w(w113_27),.acc(r113_27),.res(r113_28),.clk(clk),.wout(w113_28));
	PE pe113_29(.x(x29),.w(w113_28),.acc(r113_28),.res(r113_29),.clk(clk),.wout(w113_29));
	PE pe113_30(.x(x30),.w(w113_29),.acc(r113_29),.res(r113_30),.clk(clk),.wout(w113_30));
	PE pe113_31(.x(x31),.w(w113_30),.acc(r113_30),.res(r113_31),.clk(clk),.wout(w113_31));
	PE pe113_32(.x(x32),.w(w113_31),.acc(r113_31),.res(r113_32),.clk(clk),.wout(w113_32));
	PE pe113_33(.x(x33),.w(w113_32),.acc(r113_32),.res(r113_33),.clk(clk),.wout(w113_33));
	PE pe113_34(.x(x34),.w(w113_33),.acc(r113_33),.res(r113_34),.clk(clk),.wout(w113_34));
	PE pe113_35(.x(x35),.w(w113_34),.acc(r113_34),.res(r113_35),.clk(clk),.wout(w113_35));
	PE pe113_36(.x(x36),.w(w113_35),.acc(r113_35),.res(r113_36),.clk(clk),.wout(w113_36));
	PE pe113_37(.x(x37),.w(w113_36),.acc(r113_36),.res(r113_37),.clk(clk),.wout(w113_37));
	PE pe113_38(.x(x38),.w(w113_37),.acc(r113_37),.res(r113_38),.clk(clk),.wout(w113_38));
	PE pe113_39(.x(x39),.w(w113_38),.acc(r113_38),.res(r113_39),.clk(clk),.wout(w113_39));
	PE pe113_40(.x(x40),.w(w113_39),.acc(r113_39),.res(r113_40),.clk(clk),.wout(w113_40));
	PE pe113_41(.x(x41),.w(w113_40),.acc(r113_40),.res(r113_41),.clk(clk),.wout(w113_41));
	PE pe113_42(.x(x42),.w(w113_41),.acc(r113_41),.res(r113_42),.clk(clk),.wout(w113_42));
	PE pe113_43(.x(x43),.w(w113_42),.acc(r113_42),.res(r113_43),.clk(clk),.wout(w113_43));
	PE pe113_44(.x(x44),.w(w113_43),.acc(r113_43),.res(r113_44),.clk(clk),.wout(w113_44));
	PE pe113_45(.x(x45),.w(w113_44),.acc(r113_44),.res(r113_45),.clk(clk),.wout(w113_45));
	PE pe113_46(.x(x46),.w(w113_45),.acc(r113_45),.res(r113_46),.clk(clk),.wout(w113_46));
	PE pe113_47(.x(x47),.w(w113_46),.acc(r113_46),.res(r113_47),.clk(clk),.wout(w113_47));
	PE pe113_48(.x(x48),.w(w113_47),.acc(r113_47),.res(r113_48),.clk(clk),.wout(w113_48));
	PE pe113_49(.x(x49),.w(w113_48),.acc(r113_48),.res(r113_49),.clk(clk),.wout(w113_49));
	PE pe113_50(.x(x50),.w(w113_49),.acc(r113_49),.res(r113_50),.clk(clk),.wout(w113_50));
	PE pe113_51(.x(x51),.w(w113_50),.acc(r113_50),.res(r113_51),.clk(clk),.wout(w113_51));
	PE pe113_52(.x(x52),.w(w113_51),.acc(r113_51),.res(r113_52),.clk(clk),.wout(w113_52));
	PE pe113_53(.x(x53),.w(w113_52),.acc(r113_52),.res(r113_53),.clk(clk),.wout(w113_53));
	PE pe113_54(.x(x54),.w(w113_53),.acc(r113_53),.res(r113_54),.clk(clk),.wout(w113_54));
	PE pe113_55(.x(x55),.w(w113_54),.acc(r113_54),.res(r113_55),.clk(clk),.wout(w113_55));
	PE pe113_56(.x(x56),.w(w113_55),.acc(r113_55),.res(r113_56),.clk(clk),.wout(w113_56));
	PE pe113_57(.x(x57),.w(w113_56),.acc(r113_56),.res(r113_57),.clk(clk),.wout(w113_57));
	PE pe113_58(.x(x58),.w(w113_57),.acc(r113_57),.res(r113_58),.clk(clk),.wout(w113_58));
	PE pe113_59(.x(x59),.w(w113_58),.acc(r113_58),.res(r113_59),.clk(clk),.wout(w113_59));
	PE pe113_60(.x(x60),.w(w113_59),.acc(r113_59),.res(r113_60),.clk(clk),.wout(w113_60));
	PE pe113_61(.x(x61),.w(w113_60),.acc(r113_60),.res(r113_61),.clk(clk),.wout(w113_61));
	PE pe113_62(.x(x62),.w(w113_61),.acc(r113_61),.res(r113_62),.clk(clk),.wout(w113_62));
	PE pe113_63(.x(x63),.w(w113_62),.acc(r113_62),.res(r113_63),.clk(clk),.wout(w113_63));
	PE pe113_64(.x(x64),.w(w113_63),.acc(r113_63),.res(r113_64),.clk(clk),.wout(w113_64));
	PE pe113_65(.x(x65),.w(w113_64),.acc(r113_64),.res(r113_65),.clk(clk),.wout(w113_65));
	PE pe113_66(.x(x66),.w(w113_65),.acc(r113_65),.res(r113_66),.clk(clk),.wout(w113_66));
	PE pe113_67(.x(x67),.w(w113_66),.acc(r113_66),.res(r113_67),.clk(clk),.wout(w113_67));
	PE pe113_68(.x(x68),.w(w113_67),.acc(r113_67),.res(r113_68),.clk(clk),.wout(w113_68));
	PE pe113_69(.x(x69),.w(w113_68),.acc(r113_68),.res(r113_69),.clk(clk),.wout(w113_69));
	PE pe113_70(.x(x70),.w(w113_69),.acc(r113_69),.res(r113_70),.clk(clk),.wout(w113_70));
	PE pe113_71(.x(x71),.w(w113_70),.acc(r113_70),.res(r113_71),.clk(clk),.wout(w113_71));
	PE pe113_72(.x(x72),.w(w113_71),.acc(r113_71),.res(r113_72),.clk(clk),.wout(w113_72));
	PE pe113_73(.x(x73),.w(w113_72),.acc(r113_72),.res(r113_73),.clk(clk),.wout(w113_73));
	PE pe113_74(.x(x74),.w(w113_73),.acc(r113_73),.res(r113_74),.clk(clk),.wout(w113_74));
	PE pe113_75(.x(x75),.w(w113_74),.acc(r113_74),.res(r113_75),.clk(clk),.wout(w113_75));
	PE pe113_76(.x(x76),.w(w113_75),.acc(r113_75),.res(r113_76),.clk(clk),.wout(w113_76));
	PE pe113_77(.x(x77),.w(w113_76),.acc(r113_76),.res(r113_77),.clk(clk),.wout(w113_77));
	PE pe113_78(.x(x78),.w(w113_77),.acc(r113_77),.res(r113_78),.clk(clk),.wout(w113_78));
	PE pe113_79(.x(x79),.w(w113_78),.acc(r113_78),.res(r113_79),.clk(clk),.wout(w113_79));
	PE pe113_80(.x(x80),.w(w113_79),.acc(r113_79),.res(r113_80),.clk(clk),.wout(w113_80));
	PE pe113_81(.x(x81),.w(w113_80),.acc(r113_80),.res(r113_81),.clk(clk),.wout(w113_81));
	PE pe113_82(.x(x82),.w(w113_81),.acc(r113_81),.res(r113_82),.clk(clk),.wout(w113_82));
	PE pe113_83(.x(x83),.w(w113_82),.acc(r113_82),.res(r113_83),.clk(clk),.wout(w113_83));
	PE pe113_84(.x(x84),.w(w113_83),.acc(r113_83),.res(r113_84),.clk(clk),.wout(w113_84));
	PE pe113_85(.x(x85),.w(w113_84),.acc(r113_84),.res(r113_85),.clk(clk),.wout(w113_85));
	PE pe113_86(.x(x86),.w(w113_85),.acc(r113_85),.res(r113_86),.clk(clk),.wout(w113_86));
	PE pe113_87(.x(x87),.w(w113_86),.acc(r113_86),.res(r113_87),.clk(clk),.wout(w113_87));
	PE pe113_88(.x(x88),.w(w113_87),.acc(r113_87),.res(r113_88),.clk(clk),.wout(w113_88));
	PE pe113_89(.x(x89),.w(w113_88),.acc(r113_88),.res(r113_89),.clk(clk),.wout(w113_89));
	PE pe113_90(.x(x90),.w(w113_89),.acc(r113_89),.res(r113_90),.clk(clk),.wout(w113_90));
	PE pe113_91(.x(x91),.w(w113_90),.acc(r113_90),.res(r113_91),.clk(clk),.wout(w113_91));
	PE pe113_92(.x(x92),.w(w113_91),.acc(r113_91),.res(r113_92),.clk(clk),.wout(w113_92));
	PE pe113_93(.x(x93),.w(w113_92),.acc(r113_92),.res(r113_93),.clk(clk),.wout(w113_93));
	PE pe113_94(.x(x94),.w(w113_93),.acc(r113_93),.res(r113_94),.clk(clk),.wout(w113_94));
	PE pe113_95(.x(x95),.w(w113_94),.acc(r113_94),.res(r113_95),.clk(clk),.wout(w113_95));
	PE pe113_96(.x(x96),.w(w113_95),.acc(r113_95),.res(r113_96),.clk(clk),.wout(w113_96));
	PE pe113_97(.x(x97),.w(w113_96),.acc(r113_96),.res(r113_97),.clk(clk),.wout(w113_97));
	PE pe113_98(.x(x98),.w(w113_97),.acc(r113_97),.res(r113_98),.clk(clk),.wout(w113_98));
	PE pe113_99(.x(x99),.w(w113_98),.acc(r113_98),.res(r113_99),.clk(clk),.wout(w113_99));
	PE pe113_100(.x(x100),.w(w113_99),.acc(r113_99),.res(r113_100),.clk(clk),.wout(w113_100));
	PE pe113_101(.x(x101),.w(w113_100),.acc(r113_100),.res(r113_101),.clk(clk),.wout(w113_101));
	PE pe113_102(.x(x102),.w(w113_101),.acc(r113_101),.res(r113_102),.clk(clk),.wout(w113_102));
	PE pe113_103(.x(x103),.w(w113_102),.acc(r113_102),.res(r113_103),.clk(clk),.wout(w113_103));
	PE pe113_104(.x(x104),.w(w113_103),.acc(r113_103),.res(r113_104),.clk(clk),.wout(w113_104));
	PE pe113_105(.x(x105),.w(w113_104),.acc(r113_104),.res(r113_105),.clk(clk),.wout(w113_105));
	PE pe113_106(.x(x106),.w(w113_105),.acc(r113_105),.res(r113_106),.clk(clk),.wout(w113_106));
	PE pe113_107(.x(x107),.w(w113_106),.acc(r113_106),.res(r113_107),.clk(clk),.wout(w113_107));
	PE pe113_108(.x(x108),.w(w113_107),.acc(r113_107),.res(r113_108),.clk(clk),.wout(w113_108));
	PE pe113_109(.x(x109),.w(w113_108),.acc(r113_108),.res(r113_109),.clk(clk),.wout(w113_109));
	PE pe113_110(.x(x110),.w(w113_109),.acc(r113_109),.res(r113_110),.clk(clk),.wout(w113_110));
	PE pe113_111(.x(x111),.w(w113_110),.acc(r113_110),.res(r113_111),.clk(clk),.wout(w113_111));
	PE pe113_112(.x(x112),.w(w113_111),.acc(r113_111),.res(r113_112),.clk(clk),.wout(w113_112));
	PE pe113_113(.x(x113),.w(w113_112),.acc(r113_112),.res(r113_113),.clk(clk),.wout(w113_113));
	PE pe113_114(.x(x114),.w(w113_113),.acc(r113_113),.res(r113_114),.clk(clk),.wout(w113_114));
	PE pe113_115(.x(x115),.w(w113_114),.acc(r113_114),.res(r113_115),.clk(clk),.wout(w113_115));
	PE pe113_116(.x(x116),.w(w113_115),.acc(r113_115),.res(r113_116),.clk(clk),.wout(w113_116));
	PE pe113_117(.x(x117),.w(w113_116),.acc(r113_116),.res(r113_117),.clk(clk),.wout(w113_117));
	PE pe113_118(.x(x118),.w(w113_117),.acc(r113_117),.res(r113_118),.clk(clk),.wout(w113_118));
	PE pe113_119(.x(x119),.w(w113_118),.acc(r113_118),.res(r113_119),.clk(clk),.wout(w113_119));
	PE pe113_120(.x(x120),.w(w113_119),.acc(r113_119),.res(r113_120),.clk(clk),.wout(w113_120));
	PE pe113_121(.x(x121),.w(w113_120),.acc(r113_120),.res(r113_121),.clk(clk),.wout(w113_121));
	PE pe113_122(.x(x122),.w(w113_121),.acc(r113_121),.res(r113_122),.clk(clk),.wout(w113_122));
	PE pe113_123(.x(x123),.w(w113_122),.acc(r113_122),.res(r113_123),.clk(clk),.wout(w113_123));
	PE pe113_124(.x(x124),.w(w113_123),.acc(r113_123),.res(r113_124),.clk(clk),.wout(w113_124));
	PE pe113_125(.x(x125),.w(w113_124),.acc(r113_124),.res(r113_125),.clk(clk),.wout(w113_125));
	PE pe113_126(.x(x126),.w(w113_125),.acc(r113_125),.res(r113_126),.clk(clk),.wout(w113_126));
	PE pe113_127(.x(x127),.w(w113_126),.acc(r113_126),.res(result113),.clk(clk),.wout(weight113));

	PE pe114_0(.x(x0),.w(w114),.acc(32'h0),.res(r114_0),.clk(clk),.wout(w114_0));
	PE pe114_1(.x(x1),.w(w114_0),.acc(r114_0),.res(r114_1),.clk(clk),.wout(w114_1));
	PE pe114_2(.x(x2),.w(w114_1),.acc(r114_1),.res(r114_2),.clk(clk),.wout(w114_2));
	PE pe114_3(.x(x3),.w(w114_2),.acc(r114_2),.res(r114_3),.clk(clk),.wout(w114_3));
	PE pe114_4(.x(x4),.w(w114_3),.acc(r114_3),.res(r114_4),.clk(clk),.wout(w114_4));
	PE pe114_5(.x(x5),.w(w114_4),.acc(r114_4),.res(r114_5),.clk(clk),.wout(w114_5));
	PE pe114_6(.x(x6),.w(w114_5),.acc(r114_5),.res(r114_6),.clk(clk),.wout(w114_6));
	PE pe114_7(.x(x7),.w(w114_6),.acc(r114_6),.res(r114_7),.clk(clk),.wout(w114_7));
	PE pe114_8(.x(x8),.w(w114_7),.acc(r114_7),.res(r114_8),.clk(clk),.wout(w114_8));
	PE pe114_9(.x(x9),.w(w114_8),.acc(r114_8),.res(r114_9),.clk(clk),.wout(w114_9));
	PE pe114_10(.x(x10),.w(w114_9),.acc(r114_9),.res(r114_10),.clk(clk),.wout(w114_10));
	PE pe114_11(.x(x11),.w(w114_10),.acc(r114_10),.res(r114_11),.clk(clk),.wout(w114_11));
	PE pe114_12(.x(x12),.w(w114_11),.acc(r114_11),.res(r114_12),.clk(clk),.wout(w114_12));
	PE pe114_13(.x(x13),.w(w114_12),.acc(r114_12),.res(r114_13),.clk(clk),.wout(w114_13));
	PE pe114_14(.x(x14),.w(w114_13),.acc(r114_13),.res(r114_14),.clk(clk),.wout(w114_14));
	PE pe114_15(.x(x15),.w(w114_14),.acc(r114_14),.res(r114_15),.clk(clk),.wout(w114_15));
	PE pe114_16(.x(x16),.w(w114_15),.acc(r114_15),.res(r114_16),.clk(clk),.wout(w114_16));
	PE pe114_17(.x(x17),.w(w114_16),.acc(r114_16),.res(r114_17),.clk(clk),.wout(w114_17));
	PE pe114_18(.x(x18),.w(w114_17),.acc(r114_17),.res(r114_18),.clk(clk),.wout(w114_18));
	PE pe114_19(.x(x19),.w(w114_18),.acc(r114_18),.res(r114_19),.clk(clk),.wout(w114_19));
	PE pe114_20(.x(x20),.w(w114_19),.acc(r114_19),.res(r114_20),.clk(clk),.wout(w114_20));
	PE pe114_21(.x(x21),.w(w114_20),.acc(r114_20),.res(r114_21),.clk(clk),.wout(w114_21));
	PE pe114_22(.x(x22),.w(w114_21),.acc(r114_21),.res(r114_22),.clk(clk),.wout(w114_22));
	PE pe114_23(.x(x23),.w(w114_22),.acc(r114_22),.res(r114_23),.clk(clk),.wout(w114_23));
	PE pe114_24(.x(x24),.w(w114_23),.acc(r114_23),.res(r114_24),.clk(clk),.wout(w114_24));
	PE pe114_25(.x(x25),.w(w114_24),.acc(r114_24),.res(r114_25),.clk(clk),.wout(w114_25));
	PE pe114_26(.x(x26),.w(w114_25),.acc(r114_25),.res(r114_26),.clk(clk),.wout(w114_26));
	PE pe114_27(.x(x27),.w(w114_26),.acc(r114_26),.res(r114_27),.clk(clk),.wout(w114_27));
	PE pe114_28(.x(x28),.w(w114_27),.acc(r114_27),.res(r114_28),.clk(clk),.wout(w114_28));
	PE pe114_29(.x(x29),.w(w114_28),.acc(r114_28),.res(r114_29),.clk(clk),.wout(w114_29));
	PE pe114_30(.x(x30),.w(w114_29),.acc(r114_29),.res(r114_30),.clk(clk),.wout(w114_30));
	PE pe114_31(.x(x31),.w(w114_30),.acc(r114_30),.res(r114_31),.clk(clk),.wout(w114_31));
	PE pe114_32(.x(x32),.w(w114_31),.acc(r114_31),.res(r114_32),.clk(clk),.wout(w114_32));
	PE pe114_33(.x(x33),.w(w114_32),.acc(r114_32),.res(r114_33),.clk(clk),.wout(w114_33));
	PE pe114_34(.x(x34),.w(w114_33),.acc(r114_33),.res(r114_34),.clk(clk),.wout(w114_34));
	PE pe114_35(.x(x35),.w(w114_34),.acc(r114_34),.res(r114_35),.clk(clk),.wout(w114_35));
	PE pe114_36(.x(x36),.w(w114_35),.acc(r114_35),.res(r114_36),.clk(clk),.wout(w114_36));
	PE pe114_37(.x(x37),.w(w114_36),.acc(r114_36),.res(r114_37),.clk(clk),.wout(w114_37));
	PE pe114_38(.x(x38),.w(w114_37),.acc(r114_37),.res(r114_38),.clk(clk),.wout(w114_38));
	PE pe114_39(.x(x39),.w(w114_38),.acc(r114_38),.res(r114_39),.clk(clk),.wout(w114_39));
	PE pe114_40(.x(x40),.w(w114_39),.acc(r114_39),.res(r114_40),.clk(clk),.wout(w114_40));
	PE pe114_41(.x(x41),.w(w114_40),.acc(r114_40),.res(r114_41),.clk(clk),.wout(w114_41));
	PE pe114_42(.x(x42),.w(w114_41),.acc(r114_41),.res(r114_42),.clk(clk),.wout(w114_42));
	PE pe114_43(.x(x43),.w(w114_42),.acc(r114_42),.res(r114_43),.clk(clk),.wout(w114_43));
	PE pe114_44(.x(x44),.w(w114_43),.acc(r114_43),.res(r114_44),.clk(clk),.wout(w114_44));
	PE pe114_45(.x(x45),.w(w114_44),.acc(r114_44),.res(r114_45),.clk(clk),.wout(w114_45));
	PE pe114_46(.x(x46),.w(w114_45),.acc(r114_45),.res(r114_46),.clk(clk),.wout(w114_46));
	PE pe114_47(.x(x47),.w(w114_46),.acc(r114_46),.res(r114_47),.clk(clk),.wout(w114_47));
	PE pe114_48(.x(x48),.w(w114_47),.acc(r114_47),.res(r114_48),.clk(clk),.wout(w114_48));
	PE pe114_49(.x(x49),.w(w114_48),.acc(r114_48),.res(r114_49),.clk(clk),.wout(w114_49));
	PE pe114_50(.x(x50),.w(w114_49),.acc(r114_49),.res(r114_50),.clk(clk),.wout(w114_50));
	PE pe114_51(.x(x51),.w(w114_50),.acc(r114_50),.res(r114_51),.clk(clk),.wout(w114_51));
	PE pe114_52(.x(x52),.w(w114_51),.acc(r114_51),.res(r114_52),.clk(clk),.wout(w114_52));
	PE pe114_53(.x(x53),.w(w114_52),.acc(r114_52),.res(r114_53),.clk(clk),.wout(w114_53));
	PE pe114_54(.x(x54),.w(w114_53),.acc(r114_53),.res(r114_54),.clk(clk),.wout(w114_54));
	PE pe114_55(.x(x55),.w(w114_54),.acc(r114_54),.res(r114_55),.clk(clk),.wout(w114_55));
	PE pe114_56(.x(x56),.w(w114_55),.acc(r114_55),.res(r114_56),.clk(clk),.wout(w114_56));
	PE pe114_57(.x(x57),.w(w114_56),.acc(r114_56),.res(r114_57),.clk(clk),.wout(w114_57));
	PE pe114_58(.x(x58),.w(w114_57),.acc(r114_57),.res(r114_58),.clk(clk),.wout(w114_58));
	PE pe114_59(.x(x59),.w(w114_58),.acc(r114_58),.res(r114_59),.clk(clk),.wout(w114_59));
	PE pe114_60(.x(x60),.w(w114_59),.acc(r114_59),.res(r114_60),.clk(clk),.wout(w114_60));
	PE pe114_61(.x(x61),.w(w114_60),.acc(r114_60),.res(r114_61),.clk(clk),.wout(w114_61));
	PE pe114_62(.x(x62),.w(w114_61),.acc(r114_61),.res(r114_62),.clk(clk),.wout(w114_62));
	PE pe114_63(.x(x63),.w(w114_62),.acc(r114_62),.res(r114_63),.clk(clk),.wout(w114_63));
	PE pe114_64(.x(x64),.w(w114_63),.acc(r114_63),.res(r114_64),.clk(clk),.wout(w114_64));
	PE pe114_65(.x(x65),.w(w114_64),.acc(r114_64),.res(r114_65),.clk(clk),.wout(w114_65));
	PE pe114_66(.x(x66),.w(w114_65),.acc(r114_65),.res(r114_66),.clk(clk),.wout(w114_66));
	PE pe114_67(.x(x67),.w(w114_66),.acc(r114_66),.res(r114_67),.clk(clk),.wout(w114_67));
	PE pe114_68(.x(x68),.w(w114_67),.acc(r114_67),.res(r114_68),.clk(clk),.wout(w114_68));
	PE pe114_69(.x(x69),.w(w114_68),.acc(r114_68),.res(r114_69),.clk(clk),.wout(w114_69));
	PE pe114_70(.x(x70),.w(w114_69),.acc(r114_69),.res(r114_70),.clk(clk),.wout(w114_70));
	PE pe114_71(.x(x71),.w(w114_70),.acc(r114_70),.res(r114_71),.clk(clk),.wout(w114_71));
	PE pe114_72(.x(x72),.w(w114_71),.acc(r114_71),.res(r114_72),.clk(clk),.wout(w114_72));
	PE pe114_73(.x(x73),.w(w114_72),.acc(r114_72),.res(r114_73),.clk(clk),.wout(w114_73));
	PE pe114_74(.x(x74),.w(w114_73),.acc(r114_73),.res(r114_74),.clk(clk),.wout(w114_74));
	PE pe114_75(.x(x75),.w(w114_74),.acc(r114_74),.res(r114_75),.clk(clk),.wout(w114_75));
	PE pe114_76(.x(x76),.w(w114_75),.acc(r114_75),.res(r114_76),.clk(clk),.wout(w114_76));
	PE pe114_77(.x(x77),.w(w114_76),.acc(r114_76),.res(r114_77),.clk(clk),.wout(w114_77));
	PE pe114_78(.x(x78),.w(w114_77),.acc(r114_77),.res(r114_78),.clk(clk),.wout(w114_78));
	PE pe114_79(.x(x79),.w(w114_78),.acc(r114_78),.res(r114_79),.clk(clk),.wout(w114_79));
	PE pe114_80(.x(x80),.w(w114_79),.acc(r114_79),.res(r114_80),.clk(clk),.wout(w114_80));
	PE pe114_81(.x(x81),.w(w114_80),.acc(r114_80),.res(r114_81),.clk(clk),.wout(w114_81));
	PE pe114_82(.x(x82),.w(w114_81),.acc(r114_81),.res(r114_82),.clk(clk),.wout(w114_82));
	PE pe114_83(.x(x83),.w(w114_82),.acc(r114_82),.res(r114_83),.clk(clk),.wout(w114_83));
	PE pe114_84(.x(x84),.w(w114_83),.acc(r114_83),.res(r114_84),.clk(clk),.wout(w114_84));
	PE pe114_85(.x(x85),.w(w114_84),.acc(r114_84),.res(r114_85),.clk(clk),.wout(w114_85));
	PE pe114_86(.x(x86),.w(w114_85),.acc(r114_85),.res(r114_86),.clk(clk),.wout(w114_86));
	PE pe114_87(.x(x87),.w(w114_86),.acc(r114_86),.res(r114_87),.clk(clk),.wout(w114_87));
	PE pe114_88(.x(x88),.w(w114_87),.acc(r114_87),.res(r114_88),.clk(clk),.wout(w114_88));
	PE pe114_89(.x(x89),.w(w114_88),.acc(r114_88),.res(r114_89),.clk(clk),.wout(w114_89));
	PE pe114_90(.x(x90),.w(w114_89),.acc(r114_89),.res(r114_90),.clk(clk),.wout(w114_90));
	PE pe114_91(.x(x91),.w(w114_90),.acc(r114_90),.res(r114_91),.clk(clk),.wout(w114_91));
	PE pe114_92(.x(x92),.w(w114_91),.acc(r114_91),.res(r114_92),.clk(clk),.wout(w114_92));
	PE pe114_93(.x(x93),.w(w114_92),.acc(r114_92),.res(r114_93),.clk(clk),.wout(w114_93));
	PE pe114_94(.x(x94),.w(w114_93),.acc(r114_93),.res(r114_94),.clk(clk),.wout(w114_94));
	PE pe114_95(.x(x95),.w(w114_94),.acc(r114_94),.res(r114_95),.clk(clk),.wout(w114_95));
	PE pe114_96(.x(x96),.w(w114_95),.acc(r114_95),.res(r114_96),.clk(clk),.wout(w114_96));
	PE pe114_97(.x(x97),.w(w114_96),.acc(r114_96),.res(r114_97),.clk(clk),.wout(w114_97));
	PE pe114_98(.x(x98),.w(w114_97),.acc(r114_97),.res(r114_98),.clk(clk),.wout(w114_98));
	PE pe114_99(.x(x99),.w(w114_98),.acc(r114_98),.res(r114_99),.clk(clk),.wout(w114_99));
	PE pe114_100(.x(x100),.w(w114_99),.acc(r114_99),.res(r114_100),.clk(clk),.wout(w114_100));
	PE pe114_101(.x(x101),.w(w114_100),.acc(r114_100),.res(r114_101),.clk(clk),.wout(w114_101));
	PE pe114_102(.x(x102),.w(w114_101),.acc(r114_101),.res(r114_102),.clk(clk),.wout(w114_102));
	PE pe114_103(.x(x103),.w(w114_102),.acc(r114_102),.res(r114_103),.clk(clk),.wout(w114_103));
	PE pe114_104(.x(x104),.w(w114_103),.acc(r114_103),.res(r114_104),.clk(clk),.wout(w114_104));
	PE pe114_105(.x(x105),.w(w114_104),.acc(r114_104),.res(r114_105),.clk(clk),.wout(w114_105));
	PE pe114_106(.x(x106),.w(w114_105),.acc(r114_105),.res(r114_106),.clk(clk),.wout(w114_106));
	PE pe114_107(.x(x107),.w(w114_106),.acc(r114_106),.res(r114_107),.clk(clk),.wout(w114_107));
	PE pe114_108(.x(x108),.w(w114_107),.acc(r114_107),.res(r114_108),.clk(clk),.wout(w114_108));
	PE pe114_109(.x(x109),.w(w114_108),.acc(r114_108),.res(r114_109),.clk(clk),.wout(w114_109));
	PE pe114_110(.x(x110),.w(w114_109),.acc(r114_109),.res(r114_110),.clk(clk),.wout(w114_110));
	PE pe114_111(.x(x111),.w(w114_110),.acc(r114_110),.res(r114_111),.clk(clk),.wout(w114_111));
	PE pe114_112(.x(x112),.w(w114_111),.acc(r114_111),.res(r114_112),.clk(clk),.wout(w114_112));
	PE pe114_113(.x(x113),.w(w114_112),.acc(r114_112),.res(r114_113),.clk(clk),.wout(w114_113));
	PE pe114_114(.x(x114),.w(w114_113),.acc(r114_113),.res(r114_114),.clk(clk),.wout(w114_114));
	PE pe114_115(.x(x115),.w(w114_114),.acc(r114_114),.res(r114_115),.clk(clk),.wout(w114_115));
	PE pe114_116(.x(x116),.w(w114_115),.acc(r114_115),.res(r114_116),.clk(clk),.wout(w114_116));
	PE pe114_117(.x(x117),.w(w114_116),.acc(r114_116),.res(r114_117),.clk(clk),.wout(w114_117));
	PE pe114_118(.x(x118),.w(w114_117),.acc(r114_117),.res(r114_118),.clk(clk),.wout(w114_118));
	PE pe114_119(.x(x119),.w(w114_118),.acc(r114_118),.res(r114_119),.clk(clk),.wout(w114_119));
	PE pe114_120(.x(x120),.w(w114_119),.acc(r114_119),.res(r114_120),.clk(clk),.wout(w114_120));
	PE pe114_121(.x(x121),.w(w114_120),.acc(r114_120),.res(r114_121),.clk(clk),.wout(w114_121));
	PE pe114_122(.x(x122),.w(w114_121),.acc(r114_121),.res(r114_122),.clk(clk),.wout(w114_122));
	PE pe114_123(.x(x123),.w(w114_122),.acc(r114_122),.res(r114_123),.clk(clk),.wout(w114_123));
	PE pe114_124(.x(x124),.w(w114_123),.acc(r114_123),.res(r114_124),.clk(clk),.wout(w114_124));
	PE pe114_125(.x(x125),.w(w114_124),.acc(r114_124),.res(r114_125),.clk(clk),.wout(w114_125));
	PE pe114_126(.x(x126),.w(w114_125),.acc(r114_125),.res(r114_126),.clk(clk),.wout(w114_126));
	PE pe114_127(.x(x127),.w(w114_126),.acc(r114_126),.res(result114),.clk(clk),.wout(weight114));

	PE pe115_0(.x(x0),.w(w115),.acc(32'h0),.res(r115_0),.clk(clk),.wout(w115_0));
	PE pe115_1(.x(x1),.w(w115_0),.acc(r115_0),.res(r115_1),.clk(clk),.wout(w115_1));
	PE pe115_2(.x(x2),.w(w115_1),.acc(r115_1),.res(r115_2),.clk(clk),.wout(w115_2));
	PE pe115_3(.x(x3),.w(w115_2),.acc(r115_2),.res(r115_3),.clk(clk),.wout(w115_3));
	PE pe115_4(.x(x4),.w(w115_3),.acc(r115_3),.res(r115_4),.clk(clk),.wout(w115_4));
	PE pe115_5(.x(x5),.w(w115_4),.acc(r115_4),.res(r115_5),.clk(clk),.wout(w115_5));
	PE pe115_6(.x(x6),.w(w115_5),.acc(r115_5),.res(r115_6),.clk(clk),.wout(w115_6));
	PE pe115_7(.x(x7),.w(w115_6),.acc(r115_6),.res(r115_7),.clk(clk),.wout(w115_7));
	PE pe115_8(.x(x8),.w(w115_7),.acc(r115_7),.res(r115_8),.clk(clk),.wout(w115_8));
	PE pe115_9(.x(x9),.w(w115_8),.acc(r115_8),.res(r115_9),.clk(clk),.wout(w115_9));
	PE pe115_10(.x(x10),.w(w115_9),.acc(r115_9),.res(r115_10),.clk(clk),.wout(w115_10));
	PE pe115_11(.x(x11),.w(w115_10),.acc(r115_10),.res(r115_11),.clk(clk),.wout(w115_11));
	PE pe115_12(.x(x12),.w(w115_11),.acc(r115_11),.res(r115_12),.clk(clk),.wout(w115_12));
	PE pe115_13(.x(x13),.w(w115_12),.acc(r115_12),.res(r115_13),.clk(clk),.wout(w115_13));
	PE pe115_14(.x(x14),.w(w115_13),.acc(r115_13),.res(r115_14),.clk(clk),.wout(w115_14));
	PE pe115_15(.x(x15),.w(w115_14),.acc(r115_14),.res(r115_15),.clk(clk),.wout(w115_15));
	PE pe115_16(.x(x16),.w(w115_15),.acc(r115_15),.res(r115_16),.clk(clk),.wout(w115_16));
	PE pe115_17(.x(x17),.w(w115_16),.acc(r115_16),.res(r115_17),.clk(clk),.wout(w115_17));
	PE pe115_18(.x(x18),.w(w115_17),.acc(r115_17),.res(r115_18),.clk(clk),.wout(w115_18));
	PE pe115_19(.x(x19),.w(w115_18),.acc(r115_18),.res(r115_19),.clk(clk),.wout(w115_19));
	PE pe115_20(.x(x20),.w(w115_19),.acc(r115_19),.res(r115_20),.clk(clk),.wout(w115_20));
	PE pe115_21(.x(x21),.w(w115_20),.acc(r115_20),.res(r115_21),.clk(clk),.wout(w115_21));
	PE pe115_22(.x(x22),.w(w115_21),.acc(r115_21),.res(r115_22),.clk(clk),.wout(w115_22));
	PE pe115_23(.x(x23),.w(w115_22),.acc(r115_22),.res(r115_23),.clk(clk),.wout(w115_23));
	PE pe115_24(.x(x24),.w(w115_23),.acc(r115_23),.res(r115_24),.clk(clk),.wout(w115_24));
	PE pe115_25(.x(x25),.w(w115_24),.acc(r115_24),.res(r115_25),.clk(clk),.wout(w115_25));
	PE pe115_26(.x(x26),.w(w115_25),.acc(r115_25),.res(r115_26),.clk(clk),.wout(w115_26));
	PE pe115_27(.x(x27),.w(w115_26),.acc(r115_26),.res(r115_27),.clk(clk),.wout(w115_27));
	PE pe115_28(.x(x28),.w(w115_27),.acc(r115_27),.res(r115_28),.clk(clk),.wout(w115_28));
	PE pe115_29(.x(x29),.w(w115_28),.acc(r115_28),.res(r115_29),.clk(clk),.wout(w115_29));
	PE pe115_30(.x(x30),.w(w115_29),.acc(r115_29),.res(r115_30),.clk(clk),.wout(w115_30));
	PE pe115_31(.x(x31),.w(w115_30),.acc(r115_30),.res(r115_31),.clk(clk),.wout(w115_31));
	PE pe115_32(.x(x32),.w(w115_31),.acc(r115_31),.res(r115_32),.clk(clk),.wout(w115_32));
	PE pe115_33(.x(x33),.w(w115_32),.acc(r115_32),.res(r115_33),.clk(clk),.wout(w115_33));
	PE pe115_34(.x(x34),.w(w115_33),.acc(r115_33),.res(r115_34),.clk(clk),.wout(w115_34));
	PE pe115_35(.x(x35),.w(w115_34),.acc(r115_34),.res(r115_35),.clk(clk),.wout(w115_35));
	PE pe115_36(.x(x36),.w(w115_35),.acc(r115_35),.res(r115_36),.clk(clk),.wout(w115_36));
	PE pe115_37(.x(x37),.w(w115_36),.acc(r115_36),.res(r115_37),.clk(clk),.wout(w115_37));
	PE pe115_38(.x(x38),.w(w115_37),.acc(r115_37),.res(r115_38),.clk(clk),.wout(w115_38));
	PE pe115_39(.x(x39),.w(w115_38),.acc(r115_38),.res(r115_39),.clk(clk),.wout(w115_39));
	PE pe115_40(.x(x40),.w(w115_39),.acc(r115_39),.res(r115_40),.clk(clk),.wout(w115_40));
	PE pe115_41(.x(x41),.w(w115_40),.acc(r115_40),.res(r115_41),.clk(clk),.wout(w115_41));
	PE pe115_42(.x(x42),.w(w115_41),.acc(r115_41),.res(r115_42),.clk(clk),.wout(w115_42));
	PE pe115_43(.x(x43),.w(w115_42),.acc(r115_42),.res(r115_43),.clk(clk),.wout(w115_43));
	PE pe115_44(.x(x44),.w(w115_43),.acc(r115_43),.res(r115_44),.clk(clk),.wout(w115_44));
	PE pe115_45(.x(x45),.w(w115_44),.acc(r115_44),.res(r115_45),.clk(clk),.wout(w115_45));
	PE pe115_46(.x(x46),.w(w115_45),.acc(r115_45),.res(r115_46),.clk(clk),.wout(w115_46));
	PE pe115_47(.x(x47),.w(w115_46),.acc(r115_46),.res(r115_47),.clk(clk),.wout(w115_47));
	PE pe115_48(.x(x48),.w(w115_47),.acc(r115_47),.res(r115_48),.clk(clk),.wout(w115_48));
	PE pe115_49(.x(x49),.w(w115_48),.acc(r115_48),.res(r115_49),.clk(clk),.wout(w115_49));
	PE pe115_50(.x(x50),.w(w115_49),.acc(r115_49),.res(r115_50),.clk(clk),.wout(w115_50));
	PE pe115_51(.x(x51),.w(w115_50),.acc(r115_50),.res(r115_51),.clk(clk),.wout(w115_51));
	PE pe115_52(.x(x52),.w(w115_51),.acc(r115_51),.res(r115_52),.clk(clk),.wout(w115_52));
	PE pe115_53(.x(x53),.w(w115_52),.acc(r115_52),.res(r115_53),.clk(clk),.wout(w115_53));
	PE pe115_54(.x(x54),.w(w115_53),.acc(r115_53),.res(r115_54),.clk(clk),.wout(w115_54));
	PE pe115_55(.x(x55),.w(w115_54),.acc(r115_54),.res(r115_55),.clk(clk),.wout(w115_55));
	PE pe115_56(.x(x56),.w(w115_55),.acc(r115_55),.res(r115_56),.clk(clk),.wout(w115_56));
	PE pe115_57(.x(x57),.w(w115_56),.acc(r115_56),.res(r115_57),.clk(clk),.wout(w115_57));
	PE pe115_58(.x(x58),.w(w115_57),.acc(r115_57),.res(r115_58),.clk(clk),.wout(w115_58));
	PE pe115_59(.x(x59),.w(w115_58),.acc(r115_58),.res(r115_59),.clk(clk),.wout(w115_59));
	PE pe115_60(.x(x60),.w(w115_59),.acc(r115_59),.res(r115_60),.clk(clk),.wout(w115_60));
	PE pe115_61(.x(x61),.w(w115_60),.acc(r115_60),.res(r115_61),.clk(clk),.wout(w115_61));
	PE pe115_62(.x(x62),.w(w115_61),.acc(r115_61),.res(r115_62),.clk(clk),.wout(w115_62));
	PE pe115_63(.x(x63),.w(w115_62),.acc(r115_62),.res(r115_63),.clk(clk),.wout(w115_63));
	PE pe115_64(.x(x64),.w(w115_63),.acc(r115_63),.res(r115_64),.clk(clk),.wout(w115_64));
	PE pe115_65(.x(x65),.w(w115_64),.acc(r115_64),.res(r115_65),.clk(clk),.wout(w115_65));
	PE pe115_66(.x(x66),.w(w115_65),.acc(r115_65),.res(r115_66),.clk(clk),.wout(w115_66));
	PE pe115_67(.x(x67),.w(w115_66),.acc(r115_66),.res(r115_67),.clk(clk),.wout(w115_67));
	PE pe115_68(.x(x68),.w(w115_67),.acc(r115_67),.res(r115_68),.clk(clk),.wout(w115_68));
	PE pe115_69(.x(x69),.w(w115_68),.acc(r115_68),.res(r115_69),.clk(clk),.wout(w115_69));
	PE pe115_70(.x(x70),.w(w115_69),.acc(r115_69),.res(r115_70),.clk(clk),.wout(w115_70));
	PE pe115_71(.x(x71),.w(w115_70),.acc(r115_70),.res(r115_71),.clk(clk),.wout(w115_71));
	PE pe115_72(.x(x72),.w(w115_71),.acc(r115_71),.res(r115_72),.clk(clk),.wout(w115_72));
	PE pe115_73(.x(x73),.w(w115_72),.acc(r115_72),.res(r115_73),.clk(clk),.wout(w115_73));
	PE pe115_74(.x(x74),.w(w115_73),.acc(r115_73),.res(r115_74),.clk(clk),.wout(w115_74));
	PE pe115_75(.x(x75),.w(w115_74),.acc(r115_74),.res(r115_75),.clk(clk),.wout(w115_75));
	PE pe115_76(.x(x76),.w(w115_75),.acc(r115_75),.res(r115_76),.clk(clk),.wout(w115_76));
	PE pe115_77(.x(x77),.w(w115_76),.acc(r115_76),.res(r115_77),.clk(clk),.wout(w115_77));
	PE pe115_78(.x(x78),.w(w115_77),.acc(r115_77),.res(r115_78),.clk(clk),.wout(w115_78));
	PE pe115_79(.x(x79),.w(w115_78),.acc(r115_78),.res(r115_79),.clk(clk),.wout(w115_79));
	PE pe115_80(.x(x80),.w(w115_79),.acc(r115_79),.res(r115_80),.clk(clk),.wout(w115_80));
	PE pe115_81(.x(x81),.w(w115_80),.acc(r115_80),.res(r115_81),.clk(clk),.wout(w115_81));
	PE pe115_82(.x(x82),.w(w115_81),.acc(r115_81),.res(r115_82),.clk(clk),.wout(w115_82));
	PE pe115_83(.x(x83),.w(w115_82),.acc(r115_82),.res(r115_83),.clk(clk),.wout(w115_83));
	PE pe115_84(.x(x84),.w(w115_83),.acc(r115_83),.res(r115_84),.clk(clk),.wout(w115_84));
	PE pe115_85(.x(x85),.w(w115_84),.acc(r115_84),.res(r115_85),.clk(clk),.wout(w115_85));
	PE pe115_86(.x(x86),.w(w115_85),.acc(r115_85),.res(r115_86),.clk(clk),.wout(w115_86));
	PE pe115_87(.x(x87),.w(w115_86),.acc(r115_86),.res(r115_87),.clk(clk),.wout(w115_87));
	PE pe115_88(.x(x88),.w(w115_87),.acc(r115_87),.res(r115_88),.clk(clk),.wout(w115_88));
	PE pe115_89(.x(x89),.w(w115_88),.acc(r115_88),.res(r115_89),.clk(clk),.wout(w115_89));
	PE pe115_90(.x(x90),.w(w115_89),.acc(r115_89),.res(r115_90),.clk(clk),.wout(w115_90));
	PE pe115_91(.x(x91),.w(w115_90),.acc(r115_90),.res(r115_91),.clk(clk),.wout(w115_91));
	PE pe115_92(.x(x92),.w(w115_91),.acc(r115_91),.res(r115_92),.clk(clk),.wout(w115_92));
	PE pe115_93(.x(x93),.w(w115_92),.acc(r115_92),.res(r115_93),.clk(clk),.wout(w115_93));
	PE pe115_94(.x(x94),.w(w115_93),.acc(r115_93),.res(r115_94),.clk(clk),.wout(w115_94));
	PE pe115_95(.x(x95),.w(w115_94),.acc(r115_94),.res(r115_95),.clk(clk),.wout(w115_95));
	PE pe115_96(.x(x96),.w(w115_95),.acc(r115_95),.res(r115_96),.clk(clk),.wout(w115_96));
	PE pe115_97(.x(x97),.w(w115_96),.acc(r115_96),.res(r115_97),.clk(clk),.wout(w115_97));
	PE pe115_98(.x(x98),.w(w115_97),.acc(r115_97),.res(r115_98),.clk(clk),.wout(w115_98));
	PE pe115_99(.x(x99),.w(w115_98),.acc(r115_98),.res(r115_99),.clk(clk),.wout(w115_99));
	PE pe115_100(.x(x100),.w(w115_99),.acc(r115_99),.res(r115_100),.clk(clk),.wout(w115_100));
	PE pe115_101(.x(x101),.w(w115_100),.acc(r115_100),.res(r115_101),.clk(clk),.wout(w115_101));
	PE pe115_102(.x(x102),.w(w115_101),.acc(r115_101),.res(r115_102),.clk(clk),.wout(w115_102));
	PE pe115_103(.x(x103),.w(w115_102),.acc(r115_102),.res(r115_103),.clk(clk),.wout(w115_103));
	PE pe115_104(.x(x104),.w(w115_103),.acc(r115_103),.res(r115_104),.clk(clk),.wout(w115_104));
	PE pe115_105(.x(x105),.w(w115_104),.acc(r115_104),.res(r115_105),.clk(clk),.wout(w115_105));
	PE pe115_106(.x(x106),.w(w115_105),.acc(r115_105),.res(r115_106),.clk(clk),.wout(w115_106));
	PE pe115_107(.x(x107),.w(w115_106),.acc(r115_106),.res(r115_107),.clk(clk),.wout(w115_107));
	PE pe115_108(.x(x108),.w(w115_107),.acc(r115_107),.res(r115_108),.clk(clk),.wout(w115_108));
	PE pe115_109(.x(x109),.w(w115_108),.acc(r115_108),.res(r115_109),.clk(clk),.wout(w115_109));
	PE pe115_110(.x(x110),.w(w115_109),.acc(r115_109),.res(r115_110),.clk(clk),.wout(w115_110));
	PE pe115_111(.x(x111),.w(w115_110),.acc(r115_110),.res(r115_111),.clk(clk),.wout(w115_111));
	PE pe115_112(.x(x112),.w(w115_111),.acc(r115_111),.res(r115_112),.clk(clk),.wout(w115_112));
	PE pe115_113(.x(x113),.w(w115_112),.acc(r115_112),.res(r115_113),.clk(clk),.wout(w115_113));
	PE pe115_114(.x(x114),.w(w115_113),.acc(r115_113),.res(r115_114),.clk(clk),.wout(w115_114));
	PE pe115_115(.x(x115),.w(w115_114),.acc(r115_114),.res(r115_115),.clk(clk),.wout(w115_115));
	PE pe115_116(.x(x116),.w(w115_115),.acc(r115_115),.res(r115_116),.clk(clk),.wout(w115_116));
	PE pe115_117(.x(x117),.w(w115_116),.acc(r115_116),.res(r115_117),.clk(clk),.wout(w115_117));
	PE pe115_118(.x(x118),.w(w115_117),.acc(r115_117),.res(r115_118),.clk(clk),.wout(w115_118));
	PE pe115_119(.x(x119),.w(w115_118),.acc(r115_118),.res(r115_119),.clk(clk),.wout(w115_119));
	PE pe115_120(.x(x120),.w(w115_119),.acc(r115_119),.res(r115_120),.clk(clk),.wout(w115_120));
	PE pe115_121(.x(x121),.w(w115_120),.acc(r115_120),.res(r115_121),.clk(clk),.wout(w115_121));
	PE pe115_122(.x(x122),.w(w115_121),.acc(r115_121),.res(r115_122),.clk(clk),.wout(w115_122));
	PE pe115_123(.x(x123),.w(w115_122),.acc(r115_122),.res(r115_123),.clk(clk),.wout(w115_123));
	PE pe115_124(.x(x124),.w(w115_123),.acc(r115_123),.res(r115_124),.clk(clk),.wout(w115_124));
	PE pe115_125(.x(x125),.w(w115_124),.acc(r115_124),.res(r115_125),.clk(clk),.wout(w115_125));
	PE pe115_126(.x(x126),.w(w115_125),.acc(r115_125),.res(r115_126),.clk(clk),.wout(w115_126));
	PE pe115_127(.x(x127),.w(w115_126),.acc(r115_126),.res(result115),.clk(clk),.wout(weight115));

	PE pe116_0(.x(x0),.w(w116),.acc(32'h0),.res(r116_0),.clk(clk),.wout(w116_0));
	PE pe116_1(.x(x1),.w(w116_0),.acc(r116_0),.res(r116_1),.clk(clk),.wout(w116_1));
	PE pe116_2(.x(x2),.w(w116_1),.acc(r116_1),.res(r116_2),.clk(clk),.wout(w116_2));
	PE pe116_3(.x(x3),.w(w116_2),.acc(r116_2),.res(r116_3),.clk(clk),.wout(w116_3));
	PE pe116_4(.x(x4),.w(w116_3),.acc(r116_3),.res(r116_4),.clk(clk),.wout(w116_4));
	PE pe116_5(.x(x5),.w(w116_4),.acc(r116_4),.res(r116_5),.clk(clk),.wout(w116_5));
	PE pe116_6(.x(x6),.w(w116_5),.acc(r116_5),.res(r116_6),.clk(clk),.wout(w116_6));
	PE pe116_7(.x(x7),.w(w116_6),.acc(r116_6),.res(r116_7),.clk(clk),.wout(w116_7));
	PE pe116_8(.x(x8),.w(w116_7),.acc(r116_7),.res(r116_8),.clk(clk),.wout(w116_8));
	PE pe116_9(.x(x9),.w(w116_8),.acc(r116_8),.res(r116_9),.clk(clk),.wout(w116_9));
	PE pe116_10(.x(x10),.w(w116_9),.acc(r116_9),.res(r116_10),.clk(clk),.wout(w116_10));
	PE pe116_11(.x(x11),.w(w116_10),.acc(r116_10),.res(r116_11),.clk(clk),.wout(w116_11));
	PE pe116_12(.x(x12),.w(w116_11),.acc(r116_11),.res(r116_12),.clk(clk),.wout(w116_12));
	PE pe116_13(.x(x13),.w(w116_12),.acc(r116_12),.res(r116_13),.clk(clk),.wout(w116_13));
	PE pe116_14(.x(x14),.w(w116_13),.acc(r116_13),.res(r116_14),.clk(clk),.wout(w116_14));
	PE pe116_15(.x(x15),.w(w116_14),.acc(r116_14),.res(r116_15),.clk(clk),.wout(w116_15));
	PE pe116_16(.x(x16),.w(w116_15),.acc(r116_15),.res(r116_16),.clk(clk),.wout(w116_16));
	PE pe116_17(.x(x17),.w(w116_16),.acc(r116_16),.res(r116_17),.clk(clk),.wout(w116_17));
	PE pe116_18(.x(x18),.w(w116_17),.acc(r116_17),.res(r116_18),.clk(clk),.wout(w116_18));
	PE pe116_19(.x(x19),.w(w116_18),.acc(r116_18),.res(r116_19),.clk(clk),.wout(w116_19));
	PE pe116_20(.x(x20),.w(w116_19),.acc(r116_19),.res(r116_20),.clk(clk),.wout(w116_20));
	PE pe116_21(.x(x21),.w(w116_20),.acc(r116_20),.res(r116_21),.clk(clk),.wout(w116_21));
	PE pe116_22(.x(x22),.w(w116_21),.acc(r116_21),.res(r116_22),.clk(clk),.wout(w116_22));
	PE pe116_23(.x(x23),.w(w116_22),.acc(r116_22),.res(r116_23),.clk(clk),.wout(w116_23));
	PE pe116_24(.x(x24),.w(w116_23),.acc(r116_23),.res(r116_24),.clk(clk),.wout(w116_24));
	PE pe116_25(.x(x25),.w(w116_24),.acc(r116_24),.res(r116_25),.clk(clk),.wout(w116_25));
	PE pe116_26(.x(x26),.w(w116_25),.acc(r116_25),.res(r116_26),.clk(clk),.wout(w116_26));
	PE pe116_27(.x(x27),.w(w116_26),.acc(r116_26),.res(r116_27),.clk(clk),.wout(w116_27));
	PE pe116_28(.x(x28),.w(w116_27),.acc(r116_27),.res(r116_28),.clk(clk),.wout(w116_28));
	PE pe116_29(.x(x29),.w(w116_28),.acc(r116_28),.res(r116_29),.clk(clk),.wout(w116_29));
	PE pe116_30(.x(x30),.w(w116_29),.acc(r116_29),.res(r116_30),.clk(clk),.wout(w116_30));
	PE pe116_31(.x(x31),.w(w116_30),.acc(r116_30),.res(r116_31),.clk(clk),.wout(w116_31));
	PE pe116_32(.x(x32),.w(w116_31),.acc(r116_31),.res(r116_32),.clk(clk),.wout(w116_32));
	PE pe116_33(.x(x33),.w(w116_32),.acc(r116_32),.res(r116_33),.clk(clk),.wout(w116_33));
	PE pe116_34(.x(x34),.w(w116_33),.acc(r116_33),.res(r116_34),.clk(clk),.wout(w116_34));
	PE pe116_35(.x(x35),.w(w116_34),.acc(r116_34),.res(r116_35),.clk(clk),.wout(w116_35));
	PE pe116_36(.x(x36),.w(w116_35),.acc(r116_35),.res(r116_36),.clk(clk),.wout(w116_36));
	PE pe116_37(.x(x37),.w(w116_36),.acc(r116_36),.res(r116_37),.clk(clk),.wout(w116_37));
	PE pe116_38(.x(x38),.w(w116_37),.acc(r116_37),.res(r116_38),.clk(clk),.wout(w116_38));
	PE pe116_39(.x(x39),.w(w116_38),.acc(r116_38),.res(r116_39),.clk(clk),.wout(w116_39));
	PE pe116_40(.x(x40),.w(w116_39),.acc(r116_39),.res(r116_40),.clk(clk),.wout(w116_40));
	PE pe116_41(.x(x41),.w(w116_40),.acc(r116_40),.res(r116_41),.clk(clk),.wout(w116_41));
	PE pe116_42(.x(x42),.w(w116_41),.acc(r116_41),.res(r116_42),.clk(clk),.wout(w116_42));
	PE pe116_43(.x(x43),.w(w116_42),.acc(r116_42),.res(r116_43),.clk(clk),.wout(w116_43));
	PE pe116_44(.x(x44),.w(w116_43),.acc(r116_43),.res(r116_44),.clk(clk),.wout(w116_44));
	PE pe116_45(.x(x45),.w(w116_44),.acc(r116_44),.res(r116_45),.clk(clk),.wout(w116_45));
	PE pe116_46(.x(x46),.w(w116_45),.acc(r116_45),.res(r116_46),.clk(clk),.wout(w116_46));
	PE pe116_47(.x(x47),.w(w116_46),.acc(r116_46),.res(r116_47),.clk(clk),.wout(w116_47));
	PE pe116_48(.x(x48),.w(w116_47),.acc(r116_47),.res(r116_48),.clk(clk),.wout(w116_48));
	PE pe116_49(.x(x49),.w(w116_48),.acc(r116_48),.res(r116_49),.clk(clk),.wout(w116_49));
	PE pe116_50(.x(x50),.w(w116_49),.acc(r116_49),.res(r116_50),.clk(clk),.wout(w116_50));
	PE pe116_51(.x(x51),.w(w116_50),.acc(r116_50),.res(r116_51),.clk(clk),.wout(w116_51));
	PE pe116_52(.x(x52),.w(w116_51),.acc(r116_51),.res(r116_52),.clk(clk),.wout(w116_52));
	PE pe116_53(.x(x53),.w(w116_52),.acc(r116_52),.res(r116_53),.clk(clk),.wout(w116_53));
	PE pe116_54(.x(x54),.w(w116_53),.acc(r116_53),.res(r116_54),.clk(clk),.wout(w116_54));
	PE pe116_55(.x(x55),.w(w116_54),.acc(r116_54),.res(r116_55),.clk(clk),.wout(w116_55));
	PE pe116_56(.x(x56),.w(w116_55),.acc(r116_55),.res(r116_56),.clk(clk),.wout(w116_56));
	PE pe116_57(.x(x57),.w(w116_56),.acc(r116_56),.res(r116_57),.clk(clk),.wout(w116_57));
	PE pe116_58(.x(x58),.w(w116_57),.acc(r116_57),.res(r116_58),.clk(clk),.wout(w116_58));
	PE pe116_59(.x(x59),.w(w116_58),.acc(r116_58),.res(r116_59),.clk(clk),.wout(w116_59));
	PE pe116_60(.x(x60),.w(w116_59),.acc(r116_59),.res(r116_60),.clk(clk),.wout(w116_60));
	PE pe116_61(.x(x61),.w(w116_60),.acc(r116_60),.res(r116_61),.clk(clk),.wout(w116_61));
	PE pe116_62(.x(x62),.w(w116_61),.acc(r116_61),.res(r116_62),.clk(clk),.wout(w116_62));
	PE pe116_63(.x(x63),.w(w116_62),.acc(r116_62),.res(r116_63),.clk(clk),.wout(w116_63));
	PE pe116_64(.x(x64),.w(w116_63),.acc(r116_63),.res(r116_64),.clk(clk),.wout(w116_64));
	PE pe116_65(.x(x65),.w(w116_64),.acc(r116_64),.res(r116_65),.clk(clk),.wout(w116_65));
	PE pe116_66(.x(x66),.w(w116_65),.acc(r116_65),.res(r116_66),.clk(clk),.wout(w116_66));
	PE pe116_67(.x(x67),.w(w116_66),.acc(r116_66),.res(r116_67),.clk(clk),.wout(w116_67));
	PE pe116_68(.x(x68),.w(w116_67),.acc(r116_67),.res(r116_68),.clk(clk),.wout(w116_68));
	PE pe116_69(.x(x69),.w(w116_68),.acc(r116_68),.res(r116_69),.clk(clk),.wout(w116_69));
	PE pe116_70(.x(x70),.w(w116_69),.acc(r116_69),.res(r116_70),.clk(clk),.wout(w116_70));
	PE pe116_71(.x(x71),.w(w116_70),.acc(r116_70),.res(r116_71),.clk(clk),.wout(w116_71));
	PE pe116_72(.x(x72),.w(w116_71),.acc(r116_71),.res(r116_72),.clk(clk),.wout(w116_72));
	PE pe116_73(.x(x73),.w(w116_72),.acc(r116_72),.res(r116_73),.clk(clk),.wout(w116_73));
	PE pe116_74(.x(x74),.w(w116_73),.acc(r116_73),.res(r116_74),.clk(clk),.wout(w116_74));
	PE pe116_75(.x(x75),.w(w116_74),.acc(r116_74),.res(r116_75),.clk(clk),.wout(w116_75));
	PE pe116_76(.x(x76),.w(w116_75),.acc(r116_75),.res(r116_76),.clk(clk),.wout(w116_76));
	PE pe116_77(.x(x77),.w(w116_76),.acc(r116_76),.res(r116_77),.clk(clk),.wout(w116_77));
	PE pe116_78(.x(x78),.w(w116_77),.acc(r116_77),.res(r116_78),.clk(clk),.wout(w116_78));
	PE pe116_79(.x(x79),.w(w116_78),.acc(r116_78),.res(r116_79),.clk(clk),.wout(w116_79));
	PE pe116_80(.x(x80),.w(w116_79),.acc(r116_79),.res(r116_80),.clk(clk),.wout(w116_80));
	PE pe116_81(.x(x81),.w(w116_80),.acc(r116_80),.res(r116_81),.clk(clk),.wout(w116_81));
	PE pe116_82(.x(x82),.w(w116_81),.acc(r116_81),.res(r116_82),.clk(clk),.wout(w116_82));
	PE pe116_83(.x(x83),.w(w116_82),.acc(r116_82),.res(r116_83),.clk(clk),.wout(w116_83));
	PE pe116_84(.x(x84),.w(w116_83),.acc(r116_83),.res(r116_84),.clk(clk),.wout(w116_84));
	PE pe116_85(.x(x85),.w(w116_84),.acc(r116_84),.res(r116_85),.clk(clk),.wout(w116_85));
	PE pe116_86(.x(x86),.w(w116_85),.acc(r116_85),.res(r116_86),.clk(clk),.wout(w116_86));
	PE pe116_87(.x(x87),.w(w116_86),.acc(r116_86),.res(r116_87),.clk(clk),.wout(w116_87));
	PE pe116_88(.x(x88),.w(w116_87),.acc(r116_87),.res(r116_88),.clk(clk),.wout(w116_88));
	PE pe116_89(.x(x89),.w(w116_88),.acc(r116_88),.res(r116_89),.clk(clk),.wout(w116_89));
	PE pe116_90(.x(x90),.w(w116_89),.acc(r116_89),.res(r116_90),.clk(clk),.wout(w116_90));
	PE pe116_91(.x(x91),.w(w116_90),.acc(r116_90),.res(r116_91),.clk(clk),.wout(w116_91));
	PE pe116_92(.x(x92),.w(w116_91),.acc(r116_91),.res(r116_92),.clk(clk),.wout(w116_92));
	PE pe116_93(.x(x93),.w(w116_92),.acc(r116_92),.res(r116_93),.clk(clk),.wout(w116_93));
	PE pe116_94(.x(x94),.w(w116_93),.acc(r116_93),.res(r116_94),.clk(clk),.wout(w116_94));
	PE pe116_95(.x(x95),.w(w116_94),.acc(r116_94),.res(r116_95),.clk(clk),.wout(w116_95));
	PE pe116_96(.x(x96),.w(w116_95),.acc(r116_95),.res(r116_96),.clk(clk),.wout(w116_96));
	PE pe116_97(.x(x97),.w(w116_96),.acc(r116_96),.res(r116_97),.clk(clk),.wout(w116_97));
	PE pe116_98(.x(x98),.w(w116_97),.acc(r116_97),.res(r116_98),.clk(clk),.wout(w116_98));
	PE pe116_99(.x(x99),.w(w116_98),.acc(r116_98),.res(r116_99),.clk(clk),.wout(w116_99));
	PE pe116_100(.x(x100),.w(w116_99),.acc(r116_99),.res(r116_100),.clk(clk),.wout(w116_100));
	PE pe116_101(.x(x101),.w(w116_100),.acc(r116_100),.res(r116_101),.clk(clk),.wout(w116_101));
	PE pe116_102(.x(x102),.w(w116_101),.acc(r116_101),.res(r116_102),.clk(clk),.wout(w116_102));
	PE pe116_103(.x(x103),.w(w116_102),.acc(r116_102),.res(r116_103),.clk(clk),.wout(w116_103));
	PE pe116_104(.x(x104),.w(w116_103),.acc(r116_103),.res(r116_104),.clk(clk),.wout(w116_104));
	PE pe116_105(.x(x105),.w(w116_104),.acc(r116_104),.res(r116_105),.clk(clk),.wout(w116_105));
	PE pe116_106(.x(x106),.w(w116_105),.acc(r116_105),.res(r116_106),.clk(clk),.wout(w116_106));
	PE pe116_107(.x(x107),.w(w116_106),.acc(r116_106),.res(r116_107),.clk(clk),.wout(w116_107));
	PE pe116_108(.x(x108),.w(w116_107),.acc(r116_107),.res(r116_108),.clk(clk),.wout(w116_108));
	PE pe116_109(.x(x109),.w(w116_108),.acc(r116_108),.res(r116_109),.clk(clk),.wout(w116_109));
	PE pe116_110(.x(x110),.w(w116_109),.acc(r116_109),.res(r116_110),.clk(clk),.wout(w116_110));
	PE pe116_111(.x(x111),.w(w116_110),.acc(r116_110),.res(r116_111),.clk(clk),.wout(w116_111));
	PE pe116_112(.x(x112),.w(w116_111),.acc(r116_111),.res(r116_112),.clk(clk),.wout(w116_112));
	PE pe116_113(.x(x113),.w(w116_112),.acc(r116_112),.res(r116_113),.clk(clk),.wout(w116_113));
	PE pe116_114(.x(x114),.w(w116_113),.acc(r116_113),.res(r116_114),.clk(clk),.wout(w116_114));
	PE pe116_115(.x(x115),.w(w116_114),.acc(r116_114),.res(r116_115),.clk(clk),.wout(w116_115));
	PE pe116_116(.x(x116),.w(w116_115),.acc(r116_115),.res(r116_116),.clk(clk),.wout(w116_116));
	PE pe116_117(.x(x117),.w(w116_116),.acc(r116_116),.res(r116_117),.clk(clk),.wout(w116_117));
	PE pe116_118(.x(x118),.w(w116_117),.acc(r116_117),.res(r116_118),.clk(clk),.wout(w116_118));
	PE pe116_119(.x(x119),.w(w116_118),.acc(r116_118),.res(r116_119),.clk(clk),.wout(w116_119));
	PE pe116_120(.x(x120),.w(w116_119),.acc(r116_119),.res(r116_120),.clk(clk),.wout(w116_120));
	PE pe116_121(.x(x121),.w(w116_120),.acc(r116_120),.res(r116_121),.clk(clk),.wout(w116_121));
	PE pe116_122(.x(x122),.w(w116_121),.acc(r116_121),.res(r116_122),.clk(clk),.wout(w116_122));
	PE pe116_123(.x(x123),.w(w116_122),.acc(r116_122),.res(r116_123),.clk(clk),.wout(w116_123));
	PE pe116_124(.x(x124),.w(w116_123),.acc(r116_123),.res(r116_124),.clk(clk),.wout(w116_124));
	PE pe116_125(.x(x125),.w(w116_124),.acc(r116_124),.res(r116_125),.clk(clk),.wout(w116_125));
	PE pe116_126(.x(x126),.w(w116_125),.acc(r116_125),.res(r116_126),.clk(clk),.wout(w116_126));
	PE pe116_127(.x(x127),.w(w116_126),.acc(r116_126),.res(result116),.clk(clk),.wout(weight116));

	PE pe117_0(.x(x0),.w(w117),.acc(32'h0),.res(r117_0),.clk(clk),.wout(w117_0));
	PE pe117_1(.x(x1),.w(w117_0),.acc(r117_0),.res(r117_1),.clk(clk),.wout(w117_1));
	PE pe117_2(.x(x2),.w(w117_1),.acc(r117_1),.res(r117_2),.clk(clk),.wout(w117_2));
	PE pe117_3(.x(x3),.w(w117_2),.acc(r117_2),.res(r117_3),.clk(clk),.wout(w117_3));
	PE pe117_4(.x(x4),.w(w117_3),.acc(r117_3),.res(r117_4),.clk(clk),.wout(w117_4));
	PE pe117_5(.x(x5),.w(w117_4),.acc(r117_4),.res(r117_5),.clk(clk),.wout(w117_5));
	PE pe117_6(.x(x6),.w(w117_5),.acc(r117_5),.res(r117_6),.clk(clk),.wout(w117_6));
	PE pe117_7(.x(x7),.w(w117_6),.acc(r117_6),.res(r117_7),.clk(clk),.wout(w117_7));
	PE pe117_8(.x(x8),.w(w117_7),.acc(r117_7),.res(r117_8),.clk(clk),.wout(w117_8));
	PE pe117_9(.x(x9),.w(w117_8),.acc(r117_8),.res(r117_9),.clk(clk),.wout(w117_9));
	PE pe117_10(.x(x10),.w(w117_9),.acc(r117_9),.res(r117_10),.clk(clk),.wout(w117_10));
	PE pe117_11(.x(x11),.w(w117_10),.acc(r117_10),.res(r117_11),.clk(clk),.wout(w117_11));
	PE pe117_12(.x(x12),.w(w117_11),.acc(r117_11),.res(r117_12),.clk(clk),.wout(w117_12));
	PE pe117_13(.x(x13),.w(w117_12),.acc(r117_12),.res(r117_13),.clk(clk),.wout(w117_13));
	PE pe117_14(.x(x14),.w(w117_13),.acc(r117_13),.res(r117_14),.clk(clk),.wout(w117_14));
	PE pe117_15(.x(x15),.w(w117_14),.acc(r117_14),.res(r117_15),.clk(clk),.wout(w117_15));
	PE pe117_16(.x(x16),.w(w117_15),.acc(r117_15),.res(r117_16),.clk(clk),.wout(w117_16));
	PE pe117_17(.x(x17),.w(w117_16),.acc(r117_16),.res(r117_17),.clk(clk),.wout(w117_17));
	PE pe117_18(.x(x18),.w(w117_17),.acc(r117_17),.res(r117_18),.clk(clk),.wout(w117_18));
	PE pe117_19(.x(x19),.w(w117_18),.acc(r117_18),.res(r117_19),.clk(clk),.wout(w117_19));
	PE pe117_20(.x(x20),.w(w117_19),.acc(r117_19),.res(r117_20),.clk(clk),.wout(w117_20));
	PE pe117_21(.x(x21),.w(w117_20),.acc(r117_20),.res(r117_21),.clk(clk),.wout(w117_21));
	PE pe117_22(.x(x22),.w(w117_21),.acc(r117_21),.res(r117_22),.clk(clk),.wout(w117_22));
	PE pe117_23(.x(x23),.w(w117_22),.acc(r117_22),.res(r117_23),.clk(clk),.wout(w117_23));
	PE pe117_24(.x(x24),.w(w117_23),.acc(r117_23),.res(r117_24),.clk(clk),.wout(w117_24));
	PE pe117_25(.x(x25),.w(w117_24),.acc(r117_24),.res(r117_25),.clk(clk),.wout(w117_25));
	PE pe117_26(.x(x26),.w(w117_25),.acc(r117_25),.res(r117_26),.clk(clk),.wout(w117_26));
	PE pe117_27(.x(x27),.w(w117_26),.acc(r117_26),.res(r117_27),.clk(clk),.wout(w117_27));
	PE pe117_28(.x(x28),.w(w117_27),.acc(r117_27),.res(r117_28),.clk(clk),.wout(w117_28));
	PE pe117_29(.x(x29),.w(w117_28),.acc(r117_28),.res(r117_29),.clk(clk),.wout(w117_29));
	PE pe117_30(.x(x30),.w(w117_29),.acc(r117_29),.res(r117_30),.clk(clk),.wout(w117_30));
	PE pe117_31(.x(x31),.w(w117_30),.acc(r117_30),.res(r117_31),.clk(clk),.wout(w117_31));
	PE pe117_32(.x(x32),.w(w117_31),.acc(r117_31),.res(r117_32),.clk(clk),.wout(w117_32));
	PE pe117_33(.x(x33),.w(w117_32),.acc(r117_32),.res(r117_33),.clk(clk),.wout(w117_33));
	PE pe117_34(.x(x34),.w(w117_33),.acc(r117_33),.res(r117_34),.clk(clk),.wout(w117_34));
	PE pe117_35(.x(x35),.w(w117_34),.acc(r117_34),.res(r117_35),.clk(clk),.wout(w117_35));
	PE pe117_36(.x(x36),.w(w117_35),.acc(r117_35),.res(r117_36),.clk(clk),.wout(w117_36));
	PE pe117_37(.x(x37),.w(w117_36),.acc(r117_36),.res(r117_37),.clk(clk),.wout(w117_37));
	PE pe117_38(.x(x38),.w(w117_37),.acc(r117_37),.res(r117_38),.clk(clk),.wout(w117_38));
	PE pe117_39(.x(x39),.w(w117_38),.acc(r117_38),.res(r117_39),.clk(clk),.wout(w117_39));
	PE pe117_40(.x(x40),.w(w117_39),.acc(r117_39),.res(r117_40),.clk(clk),.wout(w117_40));
	PE pe117_41(.x(x41),.w(w117_40),.acc(r117_40),.res(r117_41),.clk(clk),.wout(w117_41));
	PE pe117_42(.x(x42),.w(w117_41),.acc(r117_41),.res(r117_42),.clk(clk),.wout(w117_42));
	PE pe117_43(.x(x43),.w(w117_42),.acc(r117_42),.res(r117_43),.clk(clk),.wout(w117_43));
	PE pe117_44(.x(x44),.w(w117_43),.acc(r117_43),.res(r117_44),.clk(clk),.wout(w117_44));
	PE pe117_45(.x(x45),.w(w117_44),.acc(r117_44),.res(r117_45),.clk(clk),.wout(w117_45));
	PE pe117_46(.x(x46),.w(w117_45),.acc(r117_45),.res(r117_46),.clk(clk),.wout(w117_46));
	PE pe117_47(.x(x47),.w(w117_46),.acc(r117_46),.res(r117_47),.clk(clk),.wout(w117_47));
	PE pe117_48(.x(x48),.w(w117_47),.acc(r117_47),.res(r117_48),.clk(clk),.wout(w117_48));
	PE pe117_49(.x(x49),.w(w117_48),.acc(r117_48),.res(r117_49),.clk(clk),.wout(w117_49));
	PE pe117_50(.x(x50),.w(w117_49),.acc(r117_49),.res(r117_50),.clk(clk),.wout(w117_50));
	PE pe117_51(.x(x51),.w(w117_50),.acc(r117_50),.res(r117_51),.clk(clk),.wout(w117_51));
	PE pe117_52(.x(x52),.w(w117_51),.acc(r117_51),.res(r117_52),.clk(clk),.wout(w117_52));
	PE pe117_53(.x(x53),.w(w117_52),.acc(r117_52),.res(r117_53),.clk(clk),.wout(w117_53));
	PE pe117_54(.x(x54),.w(w117_53),.acc(r117_53),.res(r117_54),.clk(clk),.wout(w117_54));
	PE pe117_55(.x(x55),.w(w117_54),.acc(r117_54),.res(r117_55),.clk(clk),.wout(w117_55));
	PE pe117_56(.x(x56),.w(w117_55),.acc(r117_55),.res(r117_56),.clk(clk),.wout(w117_56));
	PE pe117_57(.x(x57),.w(w117_56),.acc(r117_56),.res(r117_57),.clk(clk),.wout(w117_57));
	PE pe117_58(.x(x58),.w(w117_57),.acc(r117_57),.res(r117_58),.clk(clk),.wout(w117_58));
	PE pe117_59(.x(x59),.w(w117_58),.acc(r117_58),.res(r117_59),.clk(clk),.wout(w117_59));
	PE pe117_60(.x(x60),.w(w117_59),.acc(r117_59),.res(r117_60),.clk(clk),.wout(w117_60));
	PE pe117_61(.x(x61),.w(w117_60),.acc(r117_60),.res(r117_61),.clk(clk),.wout(w117_61));
	PE pe117_62(.x(x62),.w(w117_61),.acc(r117_61),.res(r117_62),.clk(clk),.wout(w117_62));
	PE pe117_63(.x(x63),.w(w117_62),.acc(r117_62),.res(r117_63),.clk(clk),.wout(w117_63));
	PE pe117_64(.x(x64),.w(w117_63),.acc(r117_63),.res(r117_64),.clk(clk),.wout(w117_64));
	PE pe117_65(.x(x65),.w(w117_64),.acc(r117_64),.res(r117_65),.clk(clk),.wout(w117_65));
	PE pe117_66(.x(x66),.w(w117_65),.acc(r117_65),.res(r117_66),.clk(clk),.wout(w117_66));
	PE pe117_67(.x(x67),.w(w117_66),.acc(r117_66),.res(r117_67),.clk(clk),.wout(w117_67));
	PE pe117_68(.x(x68),.w(w117_67),.acc(r117_67),.res(r117_68),.clk(clk),.wout(w117_68));
	PE pe117_69(.x(x69),.w(w117_68),.acc(r117_68),.res(r117_69),.clk(clk),.wout(w117_69));
	PE pe117_70(.x(x70),.w(w117_69),.acc(r117_69),.res(r117_70),.clk(clk),.wout(w117_70));
	PE pe117_71(.x(x71),.w(w117_70),.acc(r117_70),.res(r117_71),.clk(clk),.wout(w117_71));
	PE pe117_72(.x(x72),.w(w117_71),.acc(r117_71),.res(r117_72),.clk(clk),.wout(w117_72));
	PE pe117_73(.x(x73),.w(w117_72),.acc(r117_72),.res(r117_73),.clk(clk),.wout(w117_73));
	PE pe117_74(.x(x74),.w(w117_73),.acc(r117_73),.res(r117_74),.clk(clk),.wout(w117_74));
	PE pe117_75(.x(x75),.w(w117_74),.acc(r117_74),.res(r117_75),.clk(clk),.wout(w117_75));
	PE pe117_76(.x(x76),.w(w117_75),.acc(r117_75),.res(r117_76),.clk(clk),.wout(w117_76));
	PE pe117_77(.x(x77),.w(w117_76),.acc(r117_76),.res(r117_77),.clk(clk),.wout(w117_77));
	PE pe117_78(.x(x78),.w(w117_77),.acc(r117_77),.res(r117_78),.clk(clk),.wout(w117_78));
	PE pe117_79(.x(x79),.w(w117_78),.acc(r117_78),.res(r117_79),.clk(clk),.wout(w117_79));
	PE pe117_80(.x(x80),.w(w117_79),.acc(r117_79),.res(r117_80),.clk(clk),.wout(w117_80));
	PE pe117_81(.x(x81),.w(w117_80),.acc(r117_80),.res(r117_81),.clk(clk),.wout(w117_81));
	PE pe117_82(.x(x82),.w(w117_81),.acc(r117_81),.res(r117_82),.clk(clk),.wout(w117_82));
	PE pe117_83(.x(x83),.w(w117_82),.acc(r117_82),.res(r117_83),.clk(clk),.wout(w117_83));
	PE pe117_84(.x(x84),.w(w117_83),.acc(r117_83),.res(r117_84),.clk(clk),.wout(w117_84));
	PE pe117_85(.x(x85),.w(w117_84),.acc(r117_84),.res(r117_85),.clk(clk),.wout(w117_85));
	PE pe117_86(.x(x86),.w(w117_85),.acc(r117_85),.res(r117_86),.clk(clk),.wout(w117_86));
	PE pe117_87(.x(x87),.w(w117_86),.acc(r117_86),.res(r117_87),.clk(clk),.wout(w117_87));
	PE pe117_88(.x(x88),.w(w117_87),.acc(r117_87),.res(r117_88),.clk(clk),.wout(w117_88));
	PE pe117_89(.x(x89),.w(w117_88),.acc(r117_88),.res(r117_89),.clk(clk),.wout(w117_89));
	PE pe117_90(.x(x90),.w(w117_89),.acc(r117_89),.res(r117_90),.clk(clk),.wout(w117_90));
	PE pe117_91(.x(x91),.w(w117_90),.acc(r117_90),.res(r117_91),.clk(clk),.wout(w117_91));
	PE pe117_92(.x(x92),.w(w117_91),.acc(r117_91),.res(r117_92),.clk(clk),.wout(w117_92));
	PE pe117_93(.x(x93),.w(w117_92),.acc(r117_92),.res(r117_93),.clk(clk),.wout(w117_93));
	PE pe117_94(.x(x94),.w(w117_93),.acc(r117_93),.res(r117_94),.clk(clk),.wout(w117_94));
	PE pe117_95(.x(x95),.w(w117_94),.acc(r117_94),.res(r117_95),.clk(clk),.wout(w117_95));
	PE pe117_96(.x(x96),.w(w117_95),.acc(r117_95),.res(r117_96),.clk(clk),.wout(w117_96));
	PE pe117_97(.x(x97),.w(w117_96),.acc(r117_96),.res(r117_97),.clk(clk),.wout(w117_97));
	PE pe117_98(.x(x98),.w(w117_97),.acc(r117_97),.res(r117_98),.clk(clk),.wout(w117_98));
	PE pe117_99(.x(x99),.w(w117_98),.acc(r117_98),.res(r117_99),.clk(clk),.wout(w117_99));
	PE pe117_100(.x(x100),.w(w117_99),.acc(r117_99),.res(r117_100),.clk(clk),.wout(w117_100));
	PE pe117_101(.x(x101),.w(w117_100),.acc(r117_100),.res(r117_101),.clk(clk),.wout(w117_101));
	PE pe117_102(.x(x102),.w(w117_101),.acc(r117_101),.res(r117_102),.clk(clk),.wout(w117_102));
	PE pe117_103(.x(x103),.w(w117_102),.acc(r117_102),.res(r117_103),.clk(clk),.wout(w117_103));
	PE pe117_104(.x(x104),.w(w117_103),.acc(r117_103),.res(r117_104),.clk(clk),.wout(w117_104));
	PE pe117_105(.x(x105),.w(w117_104),.acc(r117_104),.res(r117_105),.clk(clk),.wout(w117_105));
	PE pe117_106(.x(x106),.w(w117_105),.acc(r117_105),.res(r117_106),.clk(clk),.wout(w117_106));
	PE pe117_107(.x(x107),.w(w117_106),.acc(r117_106),.res(r117_107),.clk(clk),.wout(w117_107));
	PE pe117_108(.x(x108),.w(w117_107),.acc(r117_107),.res(r117_108),.clk(clk),.wout(w117_108));
	PE pe117_109(.x(x109),.w(w117_108),.acc(r117_108),.res(r117_109),.clk(clk),.wout(w117_109));
	PE pe117_110(.x(x110),.w(w117_109),.acc(r117_109),.res(r117_110),.clk(clk),.wout(w117_110));
	PE pe117_111(.x(x111),.w(w117_110),.acc(r117_110),.res(r117_111),.clk(clk),.wout(w117_111));
	PE pe117_112(.x(x112),.w(w117_111),.acc(r117_111),.res(r117_112),.clk(clk),.wout(w117_112));
	PE pe117_113(.x(x113),.w(w117_112),.acc(r117_112),.res(r117_113),.clk(clk),.wout(w117_113));
	PE pe117_114(.x(x114),.w(w117_113),.acc(r117_113),.res(r117_114),.clk(clk),.wout(w117_114));
	PE pe117_115(.x(x115),.w(w117_114),.acc(r117_114),.res(r117_115),.clk(clk),.wout(w117_115));
	PE pe117_116(.x(x116),.w(w117_115),.acc(r117_115),.res(r117_116),.clk(clk),.wout(w117_116));
	PE pe117_117(.x(x117),.w(w117_116),.acc(r117_116),.res(r117_117),.clk(clk),.wout(w117_117));
	PE pe117_118(.x(x118),.w(w117_117),.acc(r117_117),.res(r117_118),.clk(clk),.wout(w117_118));
	PE pe117_119(.x(x119),.w(w117_118),.acc(r117_118),.res(r117_119),.clk(clk),.wout(w117_119));
	PE pe117_120(.x(x120),.w(w117_119),.acc(r117_119),.res(r117_120),.clk(clk),.wout(w117_120));
	PE pe117_121(.x(x121),.w(w117_120),.acc(r117_120),.res(r117_121),.clk(clk),.wout(w117_121));
	PE pe117_122(.x(x122),.w(w117_121),.acc(r117_121),.res(r117_122),.clk(clk),.wout(w117_122));
	PE pe117_123(.x(x123),.w(w117_122),.acc(r117_122),.res(r117_123),.clk(clk),.wout(w117_123));
	PE pe117_124(.x(x124),.w(w117_123),.acc(r117_123),.res(r117_124),.clk(clk),.wout(w117_124));
	PE pe117_125(.x(x125),.w(w117_124),.acc(r117_124),.res(r117_125),.clk(clk),.wout(w117_125));
	PE pe117_126(.x(x126),.w(w117_125),.acc(r117_125),.res(r117_126),.clk(clk),.wout(w117_126));
	PE pe117_127(.x(x127),.w(w117_126),.acc(r117_126),.res(result117),.clk(clk),.wout(weight117));

	PE pe118_0(.x(x0),.w(w118),.acc(32'h0),.res(r118_0),.clk(clk),.wout(w118_0));
	PE pe118_1(.x(x1),.w(w118_0),.acc(r118_0),.res(r118_1),.clk(clk),.wout(w118_1));
	PE pe118_2(.x(x2),.w(w118_1),.acc(r118_1),.res(r118_2),.clk(clk),.wout(w118_2));
	PE pe118_3(.x(x3),.w(w118_2),.acc(r118_2),.res(r118_3),.clk(clk),.wout(w118_3));
	PE pe118_4(.x(x4),.w(w118_3),.acc(r118_3),.res(r118_4),.clk(clk),.wout(w118_4));
	PE pe118_5(.x(x5),.w(w118_4),.acc(r118_4),.res(r118_5),.clk(clk),.wout(w118_5));
	PE pe118_6(.x(x6),.w(w118_5),.acc(r118_5),.res(r118_6),.clk(clk),.wout(w118_6));
	PE pe118_7(.x(x7),.w(w118_6),.acc(r118_6),.res(r118_7),.clk(clk),.wout(w118_7));
	PE pe118_8(.x(x8),.w(w118_7),.acc(r118_7),.res(r118_8),.clk(clk),.wout(w118_8));
	PE pe118_9(.x(x9),.w(w118_8),.acc(r118_8),.res(r118_9),.clk(clk),.wout(w118_9));
	PE pe118_10(.x(x10),.w(w118_9),.acc(r118_9),.res(r118_10),.clk(clk),.wout(w118_10));
	PE pe118_11(.x(x11),.w(w118_10),.acc(r118_10),.res(r118_11),.clk(clk),.wout(w118_11));
	PE pe118_12(.x(x12),.w(w118_11),.acc(r118_11),.res(r118_12),.clk(clk),.wout(w118_12));
	PE pe118_13(.x(x13),.w(w118_12),.acc(r118_12),.res(r118_13),.clk(clk),.wout(w118_13));
	PE pe118_14(.x(x14),.w(w118_13),.acc(r118_13),.res(r118_14),.clk(clk),.wout(w118_14));
	PE pe118_15(.x(x15),.w(w118_14),.acc(r118_14),.res(r118_15),.clk(clk),.wout(w118_15));
	PE pe118_16(.x(x16),.w(w118_15),.acc(r118_15),.res(r118_16),.clk(clk),.wout(w118_16));
	PE pe118_17(.x(x17),.w(w118_16),.acc(r118_16),.res(r118_17),.clk(clk),.wout(w118_17));
	PE pe118_18(.x(x18),.w(w118_17),.acc(r118_17),.res(r118_18),.clk(clk),.wout(w118_18));
	PE pe118_19(.x(x19),.w(w118_18),.acc(r118_18),.res(r118_19),.clk(clk),.wout(w118_19));
	PE pe118_20(.x(x20),.w(w118_19),.acc(r118_19),.res(r118_20),.clk(clk),.wout(w118_20));
	PE pe118_21(.x(x21),.w(w118_20),.acc(r118_20),.res(r118_21),.clk(clk),.wout(w118_21));
	PE pe118_22(.x(x22),.w(w118_21),.acc(r118_21),.res(r118_22),.clk(clk),.wout(w118_22));
	PE pe118_23(.x(x23),.w(w118_22),.acc(r118_22),.res(r118_23),.clk(clk),.wout(w118_23));
	PE pe118_24(.x(x24),.w(w118_23),.acc(r118_23),.res(r118_24),.clk(clk),.wout(w118_24));
	PE pe118_25(.x(x25),.w(w118_24),.acc(r118_24),.res(r118_25),.clk(clk),.wout(w118_25));
	PE pe118_26(.x(x26),.w(w118_25),.acc(r118_25),.res(r118_26),.clk(clk),.wout(w118_26));
	PE pe118_27(.x(x27),.w(w118_26),.acc(r118_26),.res(r118_27),.clk(clk),.wout(w118_27));
	PE pe118_28(.x(x28),.w(w118_27),.acc(r118_27),.res(r118_28),.clk(clk),.wout(w118_28));
	PE pe118_29(.x(x29),.w(w118_28),.acc(r118_28),.res(r118_29),.clk(clk),.wout(w118_29));
	PE pe118_30(.x(x30),.w(w118_29),.acc(r118_29),.res(r118_30),.clk(clk),.wout(w118_30));
	PE pe118_31(.x(x31),.w(w118_30),.acc(r118_30),.res(r118_31),.clk(clk),.wout(w118_31));
	PE pe118_32(.x(x32),.w(w118_31),.acc(r118_31),.res(r118_32),.clk(clk),.wout(w118_32));
	PE pe118_33(.x(x33),.w(w118_32),.acc(r118_32),.res(r118_33),.clk(clk),.wout(w118_33));
	PE pe118_34(.x(x34),.w(w118_33),.acc(r118_33),.res(r118_34),.clk(clk),.wout(w118_34));
	PE pe118_35(.x(x35),.w(w118_34),.acc(r118_34),.res(r118_35),.clk(clk),.wout(w118_35));
	PE pe118_36(.x(x36),.w(w118_35),.acc(r118_35),.res(r118_36),.clk(clk),.wout(w118_36));
	PE pe118_37(.x(x37),.w(w118_36),.acc(r118_36),.res(r118_37),.clk(clk),.wout(w118_37));
	PE pe118_38(.x(x38),.w(w118_37),.acc(r118_37),.res(r118_38),.clk(clk),.wout(w118_38));
	PE pe118_39(.x(x39),.w(w118_38),.acc(r118_38),.res(r118_39),.clk(clk),.wout(w118_39));
	PE pe118_40(.x(x40),.w(w118_39),.acc(r118_39),.res(r118_40),.clk(clk),.wout(w118_40));
	PE pe118_41(.x(x41),.w(w118_40),.acc(r118_40),.res(r118_41),.clk(clk),.wout(w118_41));
	PE pe118_42(.x(x42),.w(w118_41),.acc(r118_41),.res(r118_42),.clk(clk),.wout(w118_42));
	PE pe118_43(.x(x43),.w(w118_42),.acc(r118_42),.res(r118_43),.clk(clk),.wout(w118_43));
	PE pe118_44(.x(x44),.w(w118_43),.acc(r118_43),.res(r118_44),.clk(clk),.wout(w118_44));
	PE pe118_45(.x(x45),.w(w118_44),.acc(r118_44),.res(r118_45),.clk(clk),.wout(w118_45));
	PE pe118_46(.x(x46),.w(w118_45),.acc(r118_45),.res(r118_46),.clk(clk),.wout(w118_46));
	PE pe118_47(.x(x47),.w(w118_46),.acc(r118_46),.res(r118_47),.clk(clk),.wout(w118_47));
	PE pe118_48(.x(x48),.w(w118_47),.acc(r118_47),.res(r118_48),.clk(clk),.wout(w118_48));
	PE pe118_49(.x(x49),.w(w118_48),.acc(r118_48),.res(r118_49),.clk(clk),.wout(w118_49));
	PE pe118_50(.x(x50),.w(w118_49),.acc(r118_49),.res(r118_50),.clk(clk),.wout(w118_50));
	PE pe118_51(.x(x51),.w(w118_50),.acc(r118_50),.res(r118_51),.clk(clk),.wout(w118_51));
	PE pe118_52(.x(x52),.w(w118_51),.acc(r118_51),.res(r118_52),.clk(clk),.wout(w118_52));
	PE pe118_53(.x(x53),.w(w118_52),.acc(r118_52),.res(r118_53),.clk(clk),.wout(w118_53));
	PE pe118_54(.x(x54),.w(w118_53),.acc(r118_53),.res(r118_54),.clk(clk),.wout(w118_54));
	PE pe118_55(.x(x55),.w(w118_54),.acc(r118_54),.res(r118_55),.clk(clk),.wout(w118_55));
	PE pe118_56(.x(x56),.w(w118_55),.acc(r118_55),.res(r118_56),.clk(clk),.wout(w118_56));
	PE pe118_57(.x(x57),.w(w118_56),.acc(r118_56),.res(r118_57),.clk(clk),.wout(w118_57));
	PE pe118_58(.x(x58),.w(w118_57),.acc(r118_57),.res(r118_58),.clk(clk),.wout(w118_58));
	PE pe118_59(.x(x59),.w(w118_58),.acc(r118_58),.res(r118_59),.clk(clk),.wout(w118_59));
	PE pe118_60(.x(x60),.w(w118_59),.acc(r118_59),.res(r118_60),.clk(clk),.wout(w118_60));
	PE pe118_61(.x(x61),.w(w118_60),.acc(r118_60),.res(r118_61),.clk(clk),.wout(w118_61));
	PE pe118_62(.x(x62),.w(w118_61),.acc(r118_61),.res(r118_62),.clk(clk),.wout(w118_62));
	PE pe118_63(.x(x63),.w(w118_62),.acc(r118_62),.res(r118_63),.clk(clk),.wout(w118_63));
	PE pe118_64(.x(x64),.w(w118_63),.acc(r118_63),.res(r118_64),.clk(clk),.wout(w118_64));
	PE pe118_65(.x(x65),.w(w118_64),.acc(r118_64),.res(r118_65),.clk(clk),.wout(w118_65));
	PE pe118_66(.x(x66),.w(w118_65),.acc(r118_65),.res(r118_66),.clk(clk),.wout(w118_66));
	PE pe118_67(.x(x67),.w(w118_66),.acc(r118_66),.res(r118_67),.clk(clk),.wout(w118_67));
	PE pe118_68(.x(x68),.w(w118_67),.acc(r118_67),.res(r118_68),.clk(clk),.wout(w118_68));
	PE pe118_69(.x(x69),.w(w118_68),.acc(r118_68),.res(r118_69),.clk(clk),.wout(w118_69));
	PE pe118_70(.x(x70),.w(w118_69),.acc(r118_69),.res(r118_70),.clk(clk),.wout(w118_70));
	PE pe118_71(.x(x71),.w(w118_70),.acc(r118_70),.res(r118_71),.clk(clk),.wout(w118_71));
	PE pe118_72(.x(x72),.w(w118_71),.acc(r118_71),.res(r118_72),.clk(clk),.wout(w118_72));
	PE pe118_73(.x(x73),.w(w118_72),.acc(r118_72),.res(r118_73),.clk(clk),.wout(w118_73));
	PE pe118_74(.x(x74),.w(w118_73),.acc(r118_73),.res(r118_74),.clk(clk),.wout(w118_74));
	PE pe118_75(.x(x75),.w(w118_74),.acc(r118_74),.res(r118_75),.clk(clk),.wout(w118_75));
	PE pe118_76(.x(x76),.w(w118_75),.acc(r118_75),.res(r118_76),.clk(clk),.wout(w118_76));
	PE pe118_77(.x(x77),.w(w118_76),.acc(r118_76),.res(r118_77),.clk(clk),.wout(w118_77));
	PE pe118_78(.x(x78),.w(w118_77),.acc(r118_77),.res(r118_78),.clk(clk),.wout(w118_78));
	PE pe118_79(.x(x79),.w(w118_78),.acc(r118_78),.res(r118_79),.clk(clk),.wout(w118_79));
	PE pe118_80(.x(x80),.w(w118_79),.acc(r118_79),.res(r118_80),.clk(clk),.wout(w118_80));
	PE pe118_81(.x(x81),.w(w118_80),.acc(r118_80),.res(r118_81),.clk(clk),.wout(w118_81));
	PE pe118_82(.x(x82),.w(w118_81),.acc(r118_81),.res(r118_82),.clk(clk),.wout(w118_82));
	PE pe118_83(.x(x83),.w(w118_82),.acc(r118_82),.res(r118_83),.clk(clk),.wout(w118_83));
	PE pe118_84(.x(x84),.w(w118_83),.acc(r118_83),.res(r118_84),.clk(clk),.wout(w118_84));
	PE pe118_85(.x(x85),.w(w118_84),.acc(r118_84),.res(r118_85),.clk(clk),.wout(w118_85));
	PE pe118_86(.x(x86),.w(w118_85),.acc(r118_85),.res(r118_86),.clk(clk),.wout(w118_86));
	PE pe118_87(.x(x87),.w(w118_86),.acc(r118_86),.res(r118_87),.clk(clk),.wout(w118_87));
	PE pe118_88(.x(x88),.w(w118_87),.acc(r118_87),.res(r118_88),.clk(clk),.wout(w118_88));
	PE pe118_89(.x(x89),.w(w118_88),.acc(r118_88),.res(r118_89),.clk(clk),.wout(w118_89));
	PE pe118_90(.x(x90),.w(w118_89),.acc(r118_89),.res(r118_90),.clk(clk),.wout(w118_90));
	PE pe118_91(.x(x91),.w(w118_90),.acc(r118_90),.res(r118_91),.clk(clk),.wout(w118_91));
	PE pe118_92(.x(x92),.w(w118_91),.acc(r118_91),.res(r118_92),.clk(clk),.wout(w118_92));
	PE pe118_93(.x(x93),.w(w118_92),.acc(r118_92),.res(r118_93),.clk(clk),.wout(w118_93));
	PE pe118_94(.x(x94),.w(w118_93),.acc(r118_93),.res(r118_94),.clk(clk),.wout(w118_94));
	PE pe118_95(.x(x95),.w(w118_94),.acc(r118_94),.res(r118_95),.clk(clk),.wout(w118_95));
	PE pe118_96(.x(x96),.w(w118_95),.acc(r118_95),.res(r118_96),.clk(clk),.wout(w118_96));
	PE pe118_97(.x(x97),.w(w118_96),.acc(r118_96),.res(r118_97),.clk(clk),.wout(w118_97));
	PE pe118_98(.x(x98),.w(w118_97),.acc(r118_97),.res(r118_98),.clk(clk),.wout(w118_98));
	PE pe118_99(.x(x99),.w(w118_98),.acc(r118_98),.res(r118_99),.clk(clk),.wout(w118_99));
	PE pe118_100(.x(x100),.w(w118_99),.acc(r118_99),.res(r118_100),.clk(clk),.wout(w118_100));
	PE pe118_101(.x(x101),.w(w118_100),.acc(r118_100),.res(r118_101),.clk(clk),.wout(w118_101));
	PE pe118_102(.x(x102),.w(w118_101),.acc(r118_101),.res(r118_102),.clk(clk),.wout(w118_102));
	PE pe118_103(.x(x103),.w(w118_102),.acc(r118_102),.res(r118_103),.clk(clk),.wout(w118_103));
	PE pe118_104(.x(x104),.w(w118_103),.acc(r118_103),.res(r118_104),.clk(clk),.wout(w118_104));
	PE pe118_105(.x(x105),.w(w118_104),.acc(r118_104),.res(r118_105),.clk(clk),.wout(w118_105));
	PE pe118_106(.x(x106),.w(w118_105),.acc(r118_105),.res(r118_106),.clk(clk),.wout(w118_106));
	PE pe118_107(.x(x107),.w(w118_106),.acc(r118_106),.res(r118_107),.clk(clk),.wout(w118_107));
	PE pe118_108(.x(x108),.w(w118_107),.acc(r118_107),.res(r118_108),.clk(clk),.wout(w118_108));
	PE pe118_109(.x(x109),.w(w118_108),.acc(r118_108),.res(r118_109),.clk(clk),.wout(w118_109));
	PE pe118_110(.x(x110),.w(w118_109),.acc(r118_109),.res(r118_110),.clk(clk),.wout(w118_110));
	PE pe118_111(.x(x111),.w(w118_110),.acc(r118_110),.res(r118_111),.clk(clk),.wout(w118_111));
	PE pe118_112(.x(x112),.w(w118_111),.acc(r118_111),.res(r118_112),.clk(clk),.wout(w118_112));
	PE pe118_113(.x(x113),.w(w118_112),.acc(r118_112),.res(r118_113),.clk(clk),.wout(w118_113));
	PE pe118_114(.x(x114),.w(w118_113),.acc(r118_113),.res(r118_114),.clk(clk),.wout(w118_114));
	PE pe118_115(.x(x115),.w(w118_114),.acc(r118_114),.res(r118_115),.clk(clk),.wout(w118_115));
	PE pe118_116(.x(x116),.w(w118_115),.acc(r118_115),.res(r118_116),.clk(clk),.wout(w118_116));
	PE pe118_117(.x(x117),.w(w118_116),.acc(r118_116),.res(r118_117),.clk(clk),.wout(w118_117));
	PE pe118_118(.x(x118),.w(w118_117),.acc(r118_117),.res(r118_118),.clk(clk),.wout(w118_118));
	PE pe118_119(.x(x119),.w(w118_118),.acc(r118_118),.res(r118_119),.clk(clk),.wout(w118_119));
	PE pe118_120(.x(x120),.w(w118_119),.acc(r118_119),.res(r118_120),.clk(clk),.wout(w118_120));
	PE pe118_121(.x(x121),.w(w118_120),.acc(r118_120),.res(r118_121),.clk(clk),.wout(w118_121));
	PE pe118_122(.x(x122),.w(w118_121),.acc(r118_121),.res(r118_122),.clk(clk),.wout(w118_122));
	PE pe118_123(.x(x123),.w(w118_122),.acc(r118_122),.res(r118_123),.clk(clk),.wout(w118_123));
	PE pe118_124(.x(x124),.w(w118_123),.acc(r118_123),.res(r118_124),.clk(clk),.wout(w118_124));
	PE pe118_125(.x(x125),.w(w118_124),.acc(r118_124),.res(r118_125),.clk(clk),.wout(w118_125));
	PE pe118_126(.x(x126),.w(w118_125),.acc(r118_125),.res(r118_126),.clk(clk),.wout(w118_126));
	PE pe118_127(.x(x127),.w(w118_126),.acc(r118_126),.res(result118),.clk(clk),.wout(weight118));

	PE pe119_0(.x(x0),.w(w119),.acc(32'h0),.res(r119_0),.clk(clk),.wout(w119_0));
	PE pe119_1(.x(x1),.w(w119_0),.acc(r119_0),.res(r119_1),.clk(clk),.wout(w119_1));
	PE pe119_2(.x(x2),.w(w119_1),.acc(r119_1),.res(r119_2),.clk(clk),.wout(w119_2));
	PE pe119_3(.x(x3),.w(w119_2),.acc(r119_2),.res(r119_3),.clk(clk),.wout(w119_3));
	PE pe119_4(.x(x4),.w(w119_3),.acc(r119_3),.res(r119_4),.clk(clk),.wout(w119_4));
	PE pe119_5(.x(x5),.w(w119_4),.acc(r119_4),.res(r119_5),.clk(clk),.wout(w119_5));
	PE pe119_6(.x(x6),.w(w119_5),.acc(r119_5),.res(r119_6),.clk(clk),.wout(w119_6));
	PE pe119_7(.x(x7),.w(w119_6),.acc(r119_6),.res(r119_7),.clk(clk),.wout(w119_7));
	PE pe119_8(.x(x8),.w(w119_7),.acc(r119_7),.res(r119_8),.clk(clk),.wout(w119_8));
	PE pe119_9(.x(x9),.w(w119_8),.acc(r119_8),.res(r119_9),.clk(clk),.wout(w119_9));
	PE pe119_10(.x(x10),.w(w119_9),.acc(r119_9),.res(r119_10),.clk(clk),.wout(w119_10));
	PE pe119_11(.x(x11),.w(w119_10),.acc(r119_10),.res(r119_11),.clk(clk),.wout(w119_11));
	PE pe119_12(.x(x12),.w(w119_11),.acc(r119_11),.res(r119_12),.clk(clk),.wout(w119_12));
	PE pe119_13(.x(x13),.w(w119_12),.acc(r119_12),.res(r119_13),.clk(clk),.wout(w119_13));
	PE pe119_14(.x(x14),.w(w119_13),.acc(r119_13),.res(r119_14),.clk(clk),.wout(w119_14));
	PE pe119_15(.x(x15),.w(w119_14),.acc(r119_14),.res(r119_15),.clk(clk),.wout(w119_15));
	PE pe119_16(.x(x16),.w(w119_15),.acc(r119_15),.res(r119_16),.clk(clk),.wout(w119_16));
	PE pe119_17(.x(x17),.w(w119_16),.acc(r119_16),.res(r119_17),.clk(clk),.wout(w119_17));
	PE pe119_18(.x(x18),.w(w119_17),.acc(r119_17),.res(r119_18),.clk(clk),.wout(w119_18));
	PE pe119_19(.x(x19),.w(w119_18),.acc(r119_18),.res(r119_19),.clk(clk),.wout(w119_19));
	PE pe119_20(.x(x20),.w(w119_19),.acc(r119_19),.res(r119_20),.clk(clk),.wout(w119_20));
	PE pe119_21(.x(x21),.w(w119_20),.acc(r119_20),.res(r119_21),.clk(clk),.wout(w119_21));
	PE pe119_22(.x(x22),.w(w119_21),.acc(r119_21),.res(r119_22),.clk(clk),.wout(w119_22));
	PE pe119_23(.x(x23),.w(w119_22),.acc(r119_22),.res(r119_23),.clk(clk),.wout(w119_23));
	PE pe119_24(.x(x24),.w(w119_23),.acc(r119_23),.res(r119_24),.clk(clk),.wout(w119_24));
	PE pe119_25(.x(x25),.w(w119_24),.acc(r119_24),.res(r119_25),.clk(clk),.wout(w119_25));
	PE pe119_26(.x(x26),.w(w119_25),.acc(r119_25),.res(r119_26),.clk(clk),.wout(w119_26));
	PE pe119_27(.x(x27),.w(w119_26),.acc(r119_26),.res(r119_27),.clk(clk),.wout(w119_27));
	PE pe119_28(.x(x28),.w(w119_27),.acc(r119_27),.res(r119_28),.clk(clk),.wout(w119_28));
	PE pe119_29(.x(x29),.w(w119_28),.acc(r119_28),.res(r119_29),.clk(clk),.wout(w119_29));
	PE pe119_30(.x(x30),.w(w119_29),.acc(r119_29),.res(r119_30),.clk(clk),.wout(w119_30));
	PE pe119_31(.x(x31),.w(w119_30),.acc(r119_30),.res(r119_31),.clk(clk),.wout(w119_31));
	PE pe119_32(.x(x32),.w(w119_31),.acc(r119_31),.res(r119_32),.clk(clk),.wout(w119_32));
	PE pe119_33(.x(x33),.w(w119_32),.acc(r119_32),.res(r119_33),.clk(clk),.wout(w119_33));
	PE pe119_34(.x(x34),.w(w119_33),.acc(r119_33),.res(r119_34),.clk(clk),.wout(w119_34));
	PE pe119_35(.x(x35),.w(w119_34),.acc(r119_34),.res(r119_35),.clk(clk),.wout(w119_35));
	PE pe119_36(.x(x36),.w(w119_35),.acc(r119_35),.res(r119_36),.clk(clk),.wout(w119_36));
	PE pe119_37(.x(x37),.w(w119_36),.acc(r119_36),.res(r119_37),.clk(clk),.wout(w119_37));
	PE pe119_38(.x(x38),.w(w119_37),.acc(r119_37),.res(r119_38),.clk(clk),.wout(w119_38));
	PE pe119_39(.x(x39),.w(w119_38),.acc(r119_38),.res(r119_39),.clk(clk),.wout(w119_39));
	PE pe119_40(.x(x40),.w(w119_39),.acc(r119_39),.res(r119_40),.clk(clk),.wout(w119_40));
	PE pe119_41(.x(x41),.w(w119_40),.acc(r119_40),.res(r119_41),.clk(clk),.wout(w119_41));
	PE pe119_42(.x(x42),.w(w119_41),.acc(r119_41),.res(r119_42),.clk(clk),.wout(w119_42));
	PE pe119_43(.x(x43),.w(w119_42),.acc(r119_42),.res(r119_43),.clk(clk),.wout(w119_43));
	PE pe119_44(.x(x44),.w(w119_43),.acc(r119_43),.res(r119_44),.clk(clk),.wout(w119_44));
	PE pe119_45(.x(x45),.w(w119_44),.acc(r119_44),.res(r119_45),.clk(clk),.wout(w119_45));
	PE pe119_46(.x(x46),.w(w119_45),.acc(r119_45),.res(r119_46),.clk(clk),.wout(w119_46));
	PE pe119_47(.x(x47),.w(w119_46),.acc(r119_46),.res(r119_47),.clk(clk),.wout(w119_47));
	PE pe119_48(.x(x48),.w(w119_47),.acc(r119_47),.res(r119_48),.clk(clk),.wout(w119_48));
	PE pe119_49(.x(x49),.w(w119_48),.acc(r119_48),.res(r119_49),.clk(clk),.wout(w119_49));
	PE pe119_50(.x(x50),.w(w119_49),.acc(r119_49),.res(r119_50),.clk(clk),.wout(w119_50));
	PE pe119_51(.x(x51),.w(w119_50),.acc(r119_50),.res(r119_51),.clk(clk),.wout(w119_51));
	PE pe119_52(.x(x52),.w(w119_51),.acc(r119_51),.res(r119_52),.clk(clk),.wout(w119_52));
	PE pe119_53(.x(x53),.w(w119_52),.acc(r119_52),.res(r119_53),.clk(clk),.wout(w119_53));
	PE pe119_54(.x(x54),.w(w119_53),.acc(r119_53),.res(r119_54),.clk(clk),.wout(w119_54));
	PE pe119_55(.x(x55),.w(w119_54),.acc(r119_54),.res(r119_55),.clk(clk),.wout(w119_55));
	PE pe119_56(.x(x56),.w(w119_55),.acc(r119_55),.res(r119_56),.clk(clk),.wout(w119_56));
	PE pe119_57(.x(x57),.w(w119_56),.acc(r119_56),.res(r119_57),.clk(clk),.wout(w119_57));
	PE pe119_58(.x(x58),.w(w119_57),.acc(r119_57),.res(r119_58),.clk(clk),.wout(w119_58));
	PE pe119_59(.x(x59),.w(w119_58),.acc(r119_58),.res(r119_59),.clk(clk),.wout(w119_59));
	PE pe119_60(.x(x60),.w(w119_59),.acc(r119_59),.res(r119_60),.clk(clk),.wout(w119_60));
	PE pe119_61(.x(x61),.w(w119_60),.acc(r119_60),.res(r119_61),.clk(clk),.wout(w119_61));
	PE pe119_62(.x(x62),.w(w119_61),.acc(r119_61),.res(r119_62),.clk(clk),.wout(w119_62));
	PE pe119_63(.x(x63),.w(w119_62),.acc(r119_62),.res(r119_63),.clk(clk),.wout(w119_63));
	PE pe119_64(.x(x64),.w(w119_63),.acc(r119_63),.res(r119_64),.clk(clk),.wout(w119_64));
	PE pe119_65(.x(x65),.w(w119_64),.acc(r119_64),.res(r119_65),.clk(clk),.wout(w119_65));
	PE pe119_66(.x(x66),.w(w119_65),.acc(r119_65),.res(r119_66),.clk(clk),.wout(w119_66));
	PE pe119_67(.x(x67),.w(w119_66),.acc(r119_66),.res(r119_67),.clk(clk),.wout(w119_67));
	PE pe119_68(.x(x68),.w(w119_67),.acc(r119_67),.res(r119_68),.clk(clk),.wout(w119_68));
	PE pe119_69(.x(x69),.w(w119_68),.acc(r119_68),.res(r119_69),.clk(clk),.wout(w119_69));
	PE pe119_70(.x(x70),.w(w119_69),.acc(r119_69),.res(r119_70),.clk(clk),.wout(w119_70));
	PE pe119_71(.x(x71),.w(w119_70),.acc(r119_70),.res(r119_71),.clk(clk),.wout(w119_71));
	PE pe119_72(.x(x72),.w(w119_71),.acc(r119_71),.res(r119_72),.clk(clk),.wout(w119_72));
	PE pe119_73(.x(x73),.w(w119_72),.acc(r119_72),.res(r119_73),.clk(clk),.wout(w119_73));
	PE pe119_74(.x(x74),.w(w119_73),.acc(r119_73),.res(r119_74),.clk(clk),.wout(w119_74));
	PE pe119_75(.x(x75),.w(w119_74),.acc(r119_74),.res(r119_75),.clk(clk),.wout(w119_75));
	PE pe119_76(.x(x76),.w(w119_75),.acc(r119_75),.res(r119_76),.clk(clk),.wout(w119_76));
	PE pe119_77(.x(x77),.w(w119_76),.acc(r119_76),.res(r119_77),.clk(clk),.wout(w119_77));
	PE pe119_78(.x(x78),.w(w119_77),.acc(r119_77),.res(r119_78),.clk(clk),.wout(w119_78));
	PE pe119_79(.x(x79),.w(w119_78),.acc(r119_78),.res(r119_79),.clk(clk),.wout(w119_79));
	PE pe119_80(.x(x80),.w(w119_79),.acc(r119_79),.res(r119_80),.clk(clk),.wout(w119_80));
	PE pe119_81(.x(x81),.w(w119_80),.acc(r119_80),.res(r119_81),.clk(clk),.wout(w119_81));
	PE pe119_82(.x(x82),.w(w119_81),.acc(r119_81),.res(r119_82),.clk(clk),.wout(w119_82));
	PE pe119_83(.x(x83),.w(w119_82),.acc(r119_82),.res(r119_83),.clk(clk),.wout(w119_83));
	PE pe119_84(.x(x84),.w(w119_83),.acc(r119_83),.res(r119_84),.clk(clk),.wout(w119_84));
	PE pe119_85(.x(x85),.w(w119_84),.acc(r119_84),.res(r119_85),.clk(clk),.wout(w119_85));
	PE pe119_86(.x(x86),.w(w119_85),.acc(r119_85),.res(r119_86),.clk(clk),.wout(w119_86));
	PE pe119_87(.x(x87),.w(w119_86),.acc(r119_86),.res(r119_87),.clk(clk),.wout(w119_87));
	PE pe119_88(.x(x88),.w(w119_87),.acc(r119_87),.res(r119_88),.clk(clk),.wout(w119_88));
	PE pe119_89(.x(x89),.w(w119_88),.acc(r119_88),.res(r119_89),.clk(clk),.wout(w119_89));
	PE pe119_90(.x(x90),.w(w119_89),.acc(r119_89),.res(r119_90),.clk(clk),.wout(w119_90));
	PE pe119_91(.x(x91),.w(w119_90),.acc(r119_90),.res(r119_91),.clk(clk),.wout(w119_91));
	PE pe119_92(.x(x92),.w(w119_91),.acc(r119_91),.res(r119_92),.clk(clk),.wout(w119_92));
	PE pe119_93(.x(x93),.w(w119_92),.acc(r119_92),.res(r119_93),.clk(clk),.wout(w119_93));
	PE pe119_94(.x(x94),.w(w119_93),.acc(r119_93),.res(r119_94),.clk(clk),.wout(w119_94));
	PE pe119_95(.x(x95),.w(w119_94),.acc(r119_94),.res(r119_95),.clk(clk),.wout(w119_95));
	PE pe119_96(.x(x96),.w(w119_95),.acc(r119_95),.res(r119_96),.clk(clk),.wout(w119_96));
	PE pe119_97(.x(x97),.w(w119_96),.acc(r119_96),.res(r119_97),.clk(clk),.wout(w119_97));
	PE pe119_98(.x(x98),.w(w119_97),.acc(r119_97),.res(r119_98),.clk(clk),.wout(w119_98));
	PE pe119_99(.x(x99),.w(w119_98),.acc(r119_98),.res(r119_99),.clk(clk),.wout(w119_99));
	PE pe119_100(.x(x100),.w(w119_99),.acc(r119_99),.res(r119_100),.clk(clk),.wout(w119_100));
	PE pe119_101(.x(x101),.w(w119_100),.acc(r119_100),.res(r119_101),.clk(clk),.wout(w119_101));
	PE pe119_102(.x(x102),.w(w119_101),.acc(r119_101),.res(r119_102),.clk(clk),.wout(w119_102));
	PE pe119_103(.x(x103),.w(w119_102),.acc(r119_102),.res(r119_103),.clk(clk),.wout(w119_103));
	PE pe119_104(.x(x104),.w(w119_103),.acc(r119_103),.res(r119_104),.clk(clk),.wout(w119_104));
	PE pe119_105(.x(x105),.w(w119_104),.acc(r119_104),.res(r119_105),.clk(clk),.wout(w119_105));
	PE pe119_106(.x(x106),.w(w119_105),.acc(r119_105),.res(r119_106),.clk(clk),.wout(w119_106));
	PE pe119_107(.x(x107),.w(w119_106),.acc(r119_106),.res(r119_107),.clk(clk),.wout(w119_107));
	PE pe119_108(.x(x108),.w(w119_107),.acc(r119_107),.res(r119_108),.clk(clk),.wout(w119_108));
	PE pe119_109(.x(x109),.w(w119_108),.acc(r119_108),.res(r119_109),.clk(clk),.wout(w119_109));
	PE pe119_110(.x(x110),.w(w119_109),.acc(r119_109),.res(r119_110),.clk(clk),.wout(w119_110));
	PE pe119_111(.x(x111),.w(w119_110),.acc(r119_110),.res(r119_111),.clk(clk),.wout(w119_111));
	PE pe119_112(.x(x112),.w(w119_111),.acc(r119_111),.res(r119_112),.clk(clk),.wout(w119_112));
	PE pe119_113(.x(x113),.w(w119_112),.acc(r119_112),.res(r119_113),.clk(clk),.wout(w119_113));
	PE pe119_114(.x(x114),.w(w119_113),.acc(r119_113),.res(r119_114),.clk(clk),.wout(w119_114));
	PE pe119_115(.x(x115),.w(w119_114),.acc(r119_114),.res(r119_115),.clk(clk),.wout(w119_115));
	PE pe119_116(.x(x116),.w(w119_115),.acc(r119_115),.res(r119_116),.clk(clk),.wout(w119_116));
	PE pe119_117(.x(x117),.w(w119_116),.acc(r119_116),.res(r119_117),.clk(clk),.wout(w119_117));
	PE pe119_118(.x(x118),.w(w119_117),.acc(r119_117),.res(r119_118),.clk(clk),.wout(w119_118));
	PE pe119_119(.x(x119),.w(w119_118),.acc(r119_118),.res(r119_119),.clk(clk),.wout(w119_119));
	PE pe119_120(.x(x120),.w(w119_119),.acc(r119_119),.res(r119_120),.clk(clk),.wout(w119_120));
	PE pe119_121(.x(x121),.w(w119_120),.acc(r119_120),.res(r119_121),.clk(clk),.wout(w119_121));
	PE pe119_122(.x(x122),.w(w119_121),.acc(r119_121),.res(r119_122),.clk(clk),.wout(w119_122));
	PE pe119_123(.x(x123),.w(w119_122),.acc(r119_122),.res(r119_123),.clk(clk),.wout(w119_123));
	PE pe119_124(.x(x124),.w(w119_123),.acc(r119_123),.res(r119_124),.clk(clk),.wout(w119_124));
	PE pe119_125(.x(x125),.w(w119_124),.acc(r119_124),.res(r119_125),.clk(clk),.wout(w119_125));
	PE pe119_126(.x(x126),.w(w119_125),.acc(r119_125),.res(r119_126),.clk(clk),.wout(w119_126));
	PE pe119_127(.x(x127),.w(w119_126),.acc(r119_126),.res(result119),.clk(clk),.wout(weight119));

	PE pe120_0(.x(x0),.w(w120),.acc(32'h0),.res(r120_0),.clk(clk),.wout(w120_0));
	PE pe120_1(.x(x1),.w(w120_0),.acc(r120_0),.res(r120_1),.clk(clk),.wout(w120_1));
	PE pe120_2(.x(x2),.w(w120_1),.acc(r120_1),.res(r120_2),.clk(clk),.wout(w120_2));
	PE pe120_3(.x(x3),.w(w120_2),.acc(r120_2),.res(r120_3),.clk(clk),.wout(w120_3));
	PE pe120_4(.x(x4),.w(w120_3),.acc(r120_3),.res(r120_4),.clk(clk),.wout(w120_4));
	PE pe120_5(.x(x5),.w(w120_4),.acc(r120_4),.res(r120_5),.clk(clk),.wout(w120_5));
	PE pe120_6(.x(x6),.w(w120_5),.acc(r120_5),.res(r120_6),.clk(clk),.wout(w120_6));
	PE pe120_7(.x(x7),.w(w120_6),.acc(r120_6),.res(r120_7),.clk(clk),.wout(w120_7));
	PE pe120_8(.x(x8),.w(w120_7),.acc(r120_7),.res(r120_8),.clk(clk),.wout(w120_8));
	PE pe120_9(.x(x9),.w(w120_8),.acc(r120_8),.res(r120_9),.clk(clk),.wout(w120_9));
	PE pe120_10(.x(x10),.w(w120_9),.acc(r120_9),.res(r120_10),.clk(clk),.wout(w120_10));
	PE pe120_11(.x(x11),.w(w120_10),.acc(r120_10),.res(r120_11),.clk(clk),.wout(w120_11));
	PE pe120_12(.x(x12),.w(w120_11),.acc(r120_11),.res(r120_12),.clk(clk),.wout(w120_12));
	PE pe120_13(.x(x13),.w(w120_12),.acc(r120_12),.res(r120_13),.clk(clk),.wout(w120_13));
	PE pe120_14(.x(x14),.w(w120_13),.acc(r120_13),.res(r120_14),.clk(clk),.wout(w120_14));
	PE pe120_15(.x(x15),.w(w120_14),.acc(r120_14),.res(r120_15),.clk(clk),.wout(w120_15));
	PE pe120_16(.x(x16),.w(w120_15),.acc(r120_15),.res(r120_16),.clk(clk),.wout(w120_16));
	PE pe120_17(.x(x17),.w(w120_16),.acc(r120_16),.res(r120_17),.clk(clk),.wout(w120_17));
	PE pe120_18(.x(x18),.w(w120_17),.acc(r120_17),.res(r120_18),.clk(clk),.wout(w120_18));
	PE pe120_19(.x(x19),.w(w120_18),.acc(r120_18),.res(r120_19),.clk(clk),.wout(w120_19));
	PE pe120_20(.x(x20),.w(w120_19),.acc(r120_19),.res(r120_20),.clk(clk),.wout(w120_20));
	PE pe120_21(.x(x21),.w(w120_20),.acc(r120_20),.res(r120_21),.clk(clk),.wout(w120_21));
	PE pe120_22(.x(x22),.w(w120_21),.acc(r120_21),.res(r120_22),.clk(clk),.wout(w120_22));
	PE pe120_23(.x(x23),.w(w120_22),.acc(r120_22),.res(r120_23),.clk(clk),.wout(w120_23));
	PE pe120_24(.x(x24),.w(w120_23),.acc(r120_23),.res(r120_24),.clk(clk),.wout(w120_24));
	PE pe120_25(.x(x25),.w(w120_24),.acc(r120_24),.res(r120_25),.clk(clk),.wout(w120_25));
	PE pe120_26(.x(x26),.w(w120_25),.acc(r120_25),.res(r120_26),.clk(clk),.wout(w120_26));
	PE pe120_27(.x(x27),.w(w120_26),.acc(r120_26),.res(r120_27),.clk(clk),.wout(w120_27));
	PE pe120_28(.x(x28),.w(w120_27),.acc(r120_27),.res(r120_28),.clk(clk),.wout(w120_28));
	PE pe120_29(.x(x29),.w(w120_28),.acc(r120_28),.res(r120_29),.clk(clk),.wout(w120_29));
	PE pe120_30(.x(x30),.w(w120_29),.acc(r120_29),.res(r120_30),.clk(clk),.wout(w120_30));
	PE pe120_31(.x(x31),.w(w120_30),.acc(r120_30),.res(r120_31),.clk(clk),.wout(w120_31));
	PE pe120_32(.x(x32),.w(w120_31),.acc(r120_31),.res(r120_32),.clk(clk),.wout(w120_32));
	PE pe120_33(.x(x33),.w(w120_32),.acc(r120_32),.res(r120_33),.clk(clk),.wout(w120_33));
	PE pe120_34(.x(x34),.w(w120_33),.acc(r120_33),.res(r120_34),.clk(clk),.wout(w120_34));
	PE pe120_35(.x(x35),.w(w120_34),.acc(r120_34),.res(r120_35),.clk(clk),.wout(w120_35));
	PE pe120_36(.x(x36),.w(w120_35),.acc(r120_35),.res(r120_36),.clk(clk),.wout(w120_36));
	PE pe120_37(.x(x37),.w(w120_36),.acc(r120_36),.res(r120_37),.clk(clk),.wout(w120_37));
	PE pe120_38(.x(x38),.w(w120_37),.acc(r120_37),.res(r120_38),.clk(clk),.wout(w120_38));
	PE pe120_39(.x(x39),.w(w120_38),.acc(r120_38),.res(r120_39),.clk(clk),.wout(w120_39));
	PE pe120_40(.x(x40),.w(w120_39),.acc(r120_39),.res(r120_40),.clk(clk),.wout(w120_40));
	PE pe120_41(.x(x41),.w(w120_40),.acc(r120_40),.res(r120_41),.clk(clk),.wout(w120_41));
	PE pe120_42(.x(x42),.w(w120_41),.acc(r120_41),.res(r120_42),.clk(clk),.wout(w120_42));
	PE pe120_43(.x(x43),.w(w120_42),.acc(r120_42),.res(r120_43),.clk(clk),.wout(w120_43));
	PE pe120_44(.x(x44),.w(w120_43),.acc(r120_43),.res(r120_44),.clk(clk),.wout(w120_44));
	PE pe120_45(.x(x45),.w(w120_44),.acc(r120_44),.res(r120_45),.clk(clk),.wout(w120_45));
	PE pe120_46(.x(x46),.w(w120_45),.acc(r120_45),.res(r120_46),.clk(clk),.wout(w120_46));
	PE pe120_47(.x(x47),.w(w120_46),.acc(r120_46),.res(r120_47),.clk(clk),.wout(w120_47));
	PE pe120_48(.x(x48),.w(w120_47),.acc(r120_47),.res(r120_48),.clk(clk),.wout(w120_48));
	PE pe120_49(.x(x49),.w(w120_48),.acc(r120_48),.res(r120_49),.clk(clk),.wout(w120_49));
	PE pe120_50(.x(x50),.w(w120_49),.acc(r120_49),.res(r120_50),.clk(clk),.wout(w120_50));
	PE pe120_51(.x(x51),.w(w120_50),.acc(r120_50),.res(r120_51),.clk(clk),.wout(w120_51));
	PE pe120_52(.x(x52),.w(w120_51),.acc(r120_51),.res(r120_52),.clk(clk),.wout(w120_52));
	PE pe120_53(.x(x53),.w(w120_52),.acc(r120_52),.res(r120_53),.clk(clk),.wout(w120_53));
	PE pe120_54(.x(x54),.w(w120_53),.acc(r120_53),.res(r120_54),.clk(clk),.wout(w120_54));
	PE pe120_55(.x(x55),.w(w120_54),.acc(r120_54),.res(r120_55),.clk(clk),.wout(w120_55));
	PE pe120_56(.x(x56),.w(w120_55),.acc(r120_55),.res(r120_56),.clk(clk),.wout(w120_56));
	PE pe120_57(.x(x57),.w(w120_56),.acc(r120_56),.res(r120_57),.clk(clk),.wout(w120_57));
	PE pe120_58(.x(x58),.w(w120_57),.acc(r120_57),.res(r120_58),.clk(clk),.wout(w120_58));
	PE pe120_59(.x(x59),.w(w120_58),.acc(r120_58),.res(r120_59),.clk(clk),.wout(w120_59));
	PE pe120_60(.x(x60),.w(w120_59),.acc(r120_59),.res(r120_60),.clk(clk),.wout(w120_60));
	PE pe120_61(.x(x61),.w(w120_60),.acc(r120_60),.res(r120_61),.clk(clk),.wout(w120_61));
	PE pe120_62(.x(x62),.w(w120_61),.acc(r120_61),.res(r120_62),.clk(clk),.wout(w120_62));
	PE pe120_63(.x(x63),.w(w120_62),.acc(r120_62),.res(r120_63),.clk(clk),.wout(w120_63));
	PE pe120_64(.x(x64),.w(w120_63),.acc(r120_63),.res(r120_64),.clk(clk),.wout(w120_64));
	PE pe120_65(.x(x65),.w(w120_64),.acc(r120_64),.res(r120_65),.clk(clk),.wout(w120_65));
	PE pe120_66(.x(x66),.w(w120_65),.acc(r120_65),.res(r120_66),.clk(clk),.wout(w120_66));
	PE pe120_67(.x(x67),.w(w120_66),.acc(r120_66),.res(r120_67),.clk(clk),.wout(w120_67));
	PE pe120_68(.x(x68),.w(w120_67),.acc(r120_67),.res(r120_68),.clk(clk),.wout(w120_68));
	PE pe120_69(.x(x69),.w(w120_68),.acc(r120_68),.res(r120_69),.clk(clk),.wout(w120_69));
	PE pe120_70(.x(x70),.w(w120_69),.acc(r120_69),.res(r120_70),.clk(clk),.wout(w120_70));
	PE pe120_71(.x(x71),.w(w120_70),.acc(r120_70),.res(r120_71),.clk(clk),.wout(w120_71));
	PE pe120_72(.x(x72),.w(w120_71),.acc(r120_71),.res(r120_72),.clk(clk),.wout(w120_72));
	PE pe120_73(.x(x73),.w(w120_72),.acc(r120_72),.res(r120_73),.clk(clk),.wout(w120_73));
	PE pe120_74(.x(x74),.w(w120_73),.acc(r120_73),.res(r120_74),.clk(clk),.wout(w120_74));
	PE pe120_75(.x(x75),.w(w120_74),.acc(r120_74),.res(r120_75),.clk(clk),.wout(w120_75));
	PE pe120_76(.x(x76),.w(w120_75),.acc(r120_75),.res(r120_76),.clk(clk),.wout(w120_76));
	PE pe120_77(.x(x77),.w(w120_76),.acc(r120_76),.res(r120_77),.clk(clk),.wout(w120_77));
	PE pe120_78(.x(x78),.w(w120_77),.acc(r120_77),.res(r120_78),.clk(clk),.wout(w120_78));
	PE pe120_79(.x(x79),.w(w120_78),.acc(r120_78),.res(r120_79),.clk(clk),.wout(w120_79));
	PE pe120_80(.x(x80),.w(w120_79),.acc(r120_79),.res(r120_80),.clk(clk),.wout(w120_80));
	PE pe120_81(.x(x81),.w(w120_80),.acc(r120_80),.res(r120_81),.clk(clk),.wout(w120_81));
	PE pe120_82(.x(x82),.w(w120_81),.acc(r120_81),.res(r120_82),.clk(clk),.wout(w120_82));
	PE pe120_83(.x(x83),.w(w120_82),.acc(r120_82),.res(r120_83),.clk(clk),.wout(w120_83));
	PE pe120_84(.x(x84),.w(w120_83),.acc(r120_83),.res(r120_84),.clk(clk),.wout(w120_84));
	PE pe120_85(.x(x85),.w(w120_84),.acc(r120_84),.res(r120_85),.clk(clk),.wout(w120_85));
	PE pe120_86(.x(x86),.w(w120_85),.acc(r120_85),.res(r120_86),.clk(clk),.wout(w120_86));
	PE pe120_87(.x(x87),.w(w120_86),.acc(r120_86),.res(r120_87),.clk(clk),.wout(w120_87));
	PE pe120_88(.x(x88),.w(w120_87),.acc(r120_87),.res(r120_88),.clk(clk),.wout(w120_88));
	PE pe120_89(.x(x89),.w(w120_88),.acc(r120_88),.res(r120_89),.clk(clk),.wout(w120_89));
	PE pe120_90(.x(x90),.w(w120_89),.acc(r120_89),.res(r120_90),.clk(clk),.wout(w120_90));
	PE pe120_91(.x(x91),.w(w120_90),.acc(r120_90),.res(r120_91),.clk(clk),.wout(w120_91));
	PE pe120_92(.x(x92),.w(w120_91),.acc(r120_91),.res(r120_92),.clk(clk),.wout(w120_92));
	PE pe120_93(.x(x93),.w(w120_92),.acc(r120_92),.res(r120_93),.clk(clk),.wout(w120_93));
	PE pe120_94(.x(x94),.w(w120_93),.acc(r120_93),.res(r120_94),.clk(clk),.wout(w120_94));
	PE pe120_95(.x(x95),.w(w120_94),.acc(r120_94),.res(r120_95),.clk(clk),.wout(w120_95));
	PE pe120_96(.x(x96),.w(w120_95),.acc(r120_95),.res(r120_96),.clk(clk),.wout(w120_96));
	PE pe120_97(.x(x97),.w(w120_96),.acc(r120_96),.res(r120_97),.clk(clk),.wout(w120_97));
	PE pe120_98(.x(x98),.w(w120_97),.acc(r120_97),.res(r120_98),.clk(clk),.wout(w120_98));
	PE pe120_99(.x(x99),.w(w120_98),.acc(r120_98),.res(r120_99),.clk(clk),.wout(w120_99));
	PE pe120_100(.x(x100),.w(w120_99),.acc(r120_99),.res(r120_100),.clk(clk),.wout(w120_100));
	PE pe120_101(.x(x101),.w(w120_100),.acc(r120_100),.res(r120_101),.clk(clk),.wout(w120_101));
	PE pe120_102(.x(x102),.w(w120_101),.acc(r120_101),.res(r120_102),.clk(clk),.wout(w120_102));
	PE pe120_103(.x(x103),.w(w120_102),.acc(r120_102),.res(r120_103),.clk(clk),.wout(w120_103));
	PE pe120_104(.x(x104),.w(w120_103),.acc(r120_103),.res(r120_104),.clk(clk),.wout(w120_104));
	PE pe120_105(.x(x105),.w(w120_104),.acc(r120_104),.res(r120_105),.clk(clk),.wout(w120_105));
	PE pe120_106(.x(x106),.w(w120_105),.acc(r120_105),.res(r120_106),.clk(clk),.wout(w120_106));
	PE pe120_107(.x(x107),.w(w120_106),.acc(r120_106),.res(r120_107),.clk(clk),.wout(w120_107));
	PE pe120_108(.x(x108),.w(w120_107),.acc(r120_107),.res(r120_108),.clk(clk),.wout(w120_108));
	PE pe120_109(.x(x109),.w(w120_108),.acc(r120_108),.res(r120_109),.clk(clk),.wout(w120_109));
	PE pe120_110(.x(x110),.w(w120_109),.acc(r120_109),.res(r120_110),.clk(clk),.wout(w120_110));
	PE pe120_111(.x(x111),.w(w120_110),.acc(r120_110),.res(r120_111),.clk(clk),.wout(w120_111));
	PE pe120_112(.x(x112),.w(w120_111),.acc(r120_111),.res(r120_112),.clk(clk),.wout(w120_112));
	PE pe120_113(.x(x113),.w(w120_112),.acc(r120_112),.res(r120_113),.clk(clk),.wout(w120_113));
	PE pe120_114(.x(x114),.w(w120_113),.acc(r120_113),.res(r120_114),.clk(clk),.wout(w120_114));
	PE pe120_115(.x(x115),.w(w120_114),.acc(r120_114),.res(r120_115),.clk(clk),.wout(w120_115));
	PE pe120_116(.x(x116),.w(w120_115),.acc(r120_115),.res(r120_116),.clk(clk),.wout(w120_116));
	PE pe120_117(.x(x117),.w(w120_116),.acc(r120_116),.res(r120_117),.clk(clk),.wout(w120_117));
	PE pe120_118(.x(x118),.w(w120_117),.acc(r120_117),.res(r120_118),.clk(clk),.wout(w120_118));
	PE pe120_119(.x(x119),.w(w120_118),.acc(r120_118),.res(r120_119),.clk(clk),.wout(w120_119));
	PE pe120_120(.x(x120),.w(w120_119),.acc(r120_119),.res(r120_120),.clk(clk),.wout(w120_120));
	PE pe120_121(.x(x121),.w(w120_120),.acc(r120_120),.res(r120_121),.clk(clk),.wout(w120_121));
	PE pe120_122(.x(x122),.w(w120_121),.acc(r120_121),.res(r120_122),.clk(clk),.wout(w120_122));
	PE pe120_123(.x(x123),.w(w120_122),.acc(r120_122),.res(r120_123),.clk(clk),.wout(w120_123));
	PE pe120_124(.x(x124),.w(w120_123),.acc(r120_123),.res(r120_124),.clk(clk),.wout(w120_124));
	PE pe120_125(.x(x125),.w(w120_124),.acc(r120_124),.res(r120_125),.clk(clk),.wout(w120_125));
	PE pe120_126(.x(x126),.w(w120_125),.acc(r120_125),.res(r120_126),.clk(clk),.wout(w120_126));
	PE pe120_127(.x(x127),.w(w120_126),.acc(r120_126),.res(result120),.clk(clk),.wout(weight120));

	PE pe121_0(.x(x0),.w(w121),.acc(32'h0),.res(r121_0),.clk(clk),.wout(w121_0));
	PE pe121_1(.x(x1),.w(w121_0),.acc(r121_0),.res(r121_1),.clk(clk),.wout(w121_1));
	PE pe121_2(.x(x2),.w(w121_1),.acc(r121_1),.res(r121_2),.clk(clk),.wout(w121_2));
	PE pe121_3(.x(x3),.w(w121_2),.acc(r121_2),.res(r121_3),.clk(clk),.wout(w121_3));
	PE pe121_4(.x(x4),.w(w121_3),.acc(r121_3),.res(r121_4),.clk(clk),.wout(w121_4));
	PE pe121_5(.x(x5),.w(w121_4),.acc(r121_4),.res(r121_5),.clk(clk),.wout(w121_5));
	PE pe121_6(.x(x6),.w(w121_5),.acc(r121_5),.res(r121_6),.clk(clk),.wout(w121_6));
	PE pe121_7(.x(x7),.w(w121_6),.acc(r121_6),.res(r121_7),.clk(clk),.wout(w121_7));
	PE pe121_8(.x(x8),.w(w121_7),.acc(r121_7),.res(r121_8),.clk(clk),.wout(w121_8));
	PE pe121_9(.x(x9),.w(w121_8),.acc(r121_8),.res(r121_9),.clk(clk),.wout(w121_9));
	PE pe121_10(.x(x10),.w(w121_9),.acc(r121_9),.res(r121_10),.clk(clk),.wout(w121_10));
	PE pe121_11(.x(x11),.w(w121_10),.acc(r121_10),.res(r121_11),.clk(clk),.wout(w121_11));
	PE pe121_12(.x(x12),.w(w121_11),.acc(r121_11),.res(r121_12),.clk(clk),.wout(w121_12));
	PE pe121_13(.x(x13),.w(w121_12),.acc(r121_12),.res(r121_13),.clk(clk),.wout(w121_13));
	PE pe121_14(.x(x14),.w(w121_13),.acc(r121_13),.res(r121_14),.clk(clk),.wout(w121_14));
	PE pe121_15(.x(x15),.w(w121_14),.acc(r121_14),.res(r121_15),.clk(clk),.wout(w121_15));
	PE pe121_16(.x(x16),.w(w121_15),.acc(r121_15),.res(r121_16),.clk(clk),.wout(w121_16));
	PE pe121_17(.x(x17),.w(w121_16),.acc(r121_16),.res(r121_17),.clk(clk),.wout(w121_17));
	PE pe121_18(.x(x18),.w(w121_17),.acc(r121_17),.res(r121_18),.clk(clk),.wout(w121_18));
	PE pe121_19(.x(x19),.w(w121_18),.acc(r121_18),.res(r121_19),.clk(clk),.wout(w121_19));
	PE pe121_20(.x(x20),.w(w121_19),.acc(r121_19),.res(r121_20),.clk(clk),.wout(w121_20));
	PE pe121_21(.x(x21),.w(w121_20),.acc(r121_20),.res(r121_21),.clk(clk),.wout(w121_21));
	PE pe121_22(.x(x22),.w(w121_21),.acc(r121_21),.res(r121_22),.clk(clk),.wout(w121_22));
	PE pe121_23(.x(x23),.w(w121_22),.acc(r121_22),.res(r121_23),.clk(clk),.wout(w121_23));
	PE pe121_24(.x(x24),.w(w121_23),.acc(r121_23),.res(r121_24),.clk(clk),.wout(w121_24));
	PE pe121_25(.x(x25),.w(w121_24),.acc(r121_24),.res(r121_25),.clk(clk),.wout(w121_25));
	PE pe121_26(.x(x26),.w(w121_25),.acc(r121_25),.res(r121_26),.clk(clk),.wout(w121_26));
	PE pe121_27(.x(x27),.w(w121_26),.acc(r121_26),.res(r121_27),.clk(clk),.wout(w121_27));
	PE pe121_28(.x(x28),.w(w121_27),.acc(r121_27),.res(r121_28),.clk(clk),.wout(w121_28));
	PE pe121_29(.x(x29),.w(w121_28),.acc(r121_28),.res(r121_29),.clk(clk),.wout(w121_29));
	PE pe121_30(.x(x30),.w(w121_29),.acc(r121_29),.res(r121_30),.clk(clk),.wout(w121_30));
	PE pe121_31(.x(x31),.w(w121_30),.acc(r121_30),.res(r121_31),.clk(clk),.wout(w121_31));
	PE pe121_32(.x(x32),.w(w121_31),.acc(r121_31),.res(r121_32),.clk(clk),.wout(w121_32));
	PE pe121_33(.x(x33),.w(w121_32),.acc(r121_32),.res(r121_33),.clk(clk),.wout(w121_33));
	PE pe121_34(.x(x34),.w(w121_33),.acc(r121_33),.res(r121_34),.clk(clk),.wout(w121_34));
	PE pe121_35(.x(x35),.w(w121_34),.acc(r121_34),.res(r121_35),.clk(clk),.wout(w121_35));
	PE pe121_36(.x(x36),.w(w121_35),.acc(r121_35),.res(r121_36),.clk(clk),.wout(w121_36));
	PE pe121_37(.x(x37),.w(w121_36),.acc(r121_36),.res(r121_37),.clk(clk),.wout(w121_37));
	PE pe121_38(.x(x38),.w(w121_37),.acc(r121_37),.res(r121_38),.clk(clk),.wout(w121_38));
	PE pe121_39(.x(x39),.w(w121_38),.acc(r121_38),.res(r121_39),.clk(clk),.wout(w121_39));
	PE pe121_40(.x(x40),.w(w121_39),.acc(r121_39),.res(r121_40),.clk(clk),.wout(w121_40));
	PE pe121_41(.x(x41),.w(w121_40),.acc(r121_40),.res(r121_41),.clk(clk),.wout(w121_41));
	PE pe121_42(.x(x42),.w(w121_41),.acc(r121_41),.res(r121_42),.clk(clk),.wout(w121_42));
	PE pe121_43(.x(x43),.w(w121_42),.acc(r121_42),.res(r121_43),.clk(clk),.wout(w121_43));
	PE pe121_44(.x(x44),.w(w121_43),.acc(r121_43),.res(r121_44),.clk(clk),.wout(w121_44));
	PE pe121_45(.x(x45),.w(w121_44),.acc(r121_44),.res(r121_45),.clk(clk),.wout(w121_45));
	PE pe121_46(.x(x46),.w(w121_45),.acc(r121_45),.res(r121_46),.clk(clk),.wout(w121_46));
	PE pe121_47(.x(x47),.w(w121_46),.acc(r121_46),.res(r121_47),.clk(clk),.wout(w121_47));
	PE pe121_48(.x(x48),.w(w121_47),.acc(r121_47),.res(r121_48),.clk(clk),.wout(w121_48));
	PE pe121_49(.x(x49),.w(w121_48),.acc(r121_48),.res(r121_49),.clk(clk),.wout(w121_49));
	PE pe121_50(.x(x50),.w(w121_49),.acc(r121_49),.res(r121_50),.clk(clk),.wout(w121_50));
	PE pe121_51(.x(x51),.w(w121_50),.acc(r121_50),.res(r121_51),.clk(clk),.wout(w121_51));
	PE pe121_52(.x(x52),.w(w121_51),.acc(r121_51),.res(r121_52),.clk(clk),.wout(w121_52));
	PE pe121_53(.x(x53),.w(w121_52),.acc(r121_52),.res(r121_53),.clk(clk),.wout(w121_53));
	PE pe121_54(.x(x54),.w(w121_53),.acc(r121_53),.res(r121_54),.clk(clk),.wout(w121_54));
	PE pe121_55(.x(x55),.w(w121_54),.acc(r121_54),.res(r121_55),.clk(clk),.wout(w121_55));
	PE pe121_56(.x(x56),.w(w121_55),.acc(r121_55),.res(r121_56),.clk(clk),.wout(w121_56));
	PE pe121_57(.x(x57),.w(w121_56),.acc(r121_56),.res(r121_57),.clk(clk),.wout(w121_57));
	PE pe121_58(.x(x58),.w(w121_57),.acc(r121_57),.res(r121_58),.clk(clk),.wout(w121_58));
	PE pe121_59(.x(x59),.w(w121_58),.acc(r121_58),.res(r121_59),.clk(clk),.wout(w121_59));
	PE pe121_60(.x(x60),.w(w121_59),.acc(r121_59),.res(r121_60),.clk(clk),.wout(w121_60));
	PE pe121_61(.x(x61),.w(w121_60),.acc(r121_60),.res(r121_61),.clk(clk),.wout(w121_61));
	PE pe121_62(.x(x62),.w(w121_61),.acc(r121_61),.res(r121_62),.clk(clk),.wout(w121_62));
	PE pe121_63(.x(x63),.w(w121_62),.acc(r121_62),.res(r121_63),.clk(clk),.wout(w121_63));
	PE pe121_64(.x(x64),.w(w121_63),.acc(r121_63),.res(r121_64),.clk(clk),.wout(w121_64));
	PE pe121_65(.x(x65),.w(w121_64),.acc(r121_64),.res(r121_65),.clk(clk),.wout(w121_65));
	PE pe121_66(.x(x66),.w(w121_65),.acc(r121_65),.res(r121_66),.clk(clk),.wout(w121_66));
	PE pe121_67(.x(x67),.w(w121_66),.acc(r121_66),.res(r121_67),.clk(clk),.wout(w121_67));
	PE pe121_68(.x(x68),.w(w121_67),.acc(r121_67),.res(r121_68),.clk(clk),.wout(w121_68));
	PE pe121_69(.x(x69),.w(w121_68),.acc(r121_68),.res(r121_69),.clk(clk),.wout(w121_69));
	PE pe121_70(.x(x70),.w(w121_69),.acc(r121_69),.res(r121_70),.clk(clk),.wout(w121_70));
	PE pe121_71(.x(x71),.w(w121_70),.acc(r121_70),.res(r121_71),.clk(clk),.wout(w121_71));
	PE pe121_72(.x(x72),.w(w121_71),.acc(r121_71),.res(r121_72),.clk(clk),.wout(w121_72));
	PE pe121_73(.x(x73),.w(w121_72),.acc(r121_72),.res(r121_73),.clk(clk),.wout(w121_73));
	PE pe121_74(.x(x74),.w(w121_73),.acc(r121_73),.res(r121_74),.clk(clk),.wout(w121_74));
	PE pe121_75(.x(x75),.w(w121_74),.acc(r121_74),.res(r121_75),.clk(clk),.wout(w121_75));
	PE pe121_76(.x(x76),.w(w121_75),.acc(r121_75),.res(r121_76),.clk(clk),.wout(w121_76));
	PE pe121_77(.x(x77),.w(w121_76),.acc(r121_76),.res(r121_77),.clk(clk),.wout(w121_77));
	PE pe121_78(.x(x78),.w(w121_77),.acc(r121_77),.res(r121_78),.clk(clk),.wout(w121_78));
	PE pe121_79(.x(x79),.w(w121_78),.acc(r121_78),.res(r121_79),.clk(clk),.wout(w121_79));
	PE pe121_80(.x(x80),.w(w121_79),.acc(r121_79),.res(r121_80),.clk(clk),.wout(w121_80));
	PE pe121_81(.x(x81),.w(w121_80),.acc(r121_80),.res(r121_81),.clk(clk),.wout(w121_81));
	PE pe121_82(.x(x82),.w(w121_81),.acc(r121_81),.res(r121_82),.clk(clk),.wout(w121_82));
	PE pe121_83(.x(x83),.w(w121_82),.acc(r121_82),.res(r121_83),.clk(clk),.wout(w121_83));
	PE pe121_84(.x(x84),.w(w121_83),.acc(r121_83),.res(r121_84),.clk(clk),.wout(w121_84));
	PE pe121_85(.x(x85),.w(w121_84),.acc(r121_84),.res(r121_85),.clk(clk),.wout(w121_85));
	PE pe121_86(.x(x86),.w(w121_85),.acc(r121_85),.res(r121_86),.clk(clk),.wout(w121_86));
	PE pe121_87(.x(x87),.w(w121_86),.acc(r121_86),.res(r121_87),.clk(clk),.wout(w121_87));
	PE pe121_88(.x(x88),.w(w121_87),.acc(r121_87),.res(r121_88),.clk(clk),.wout(w121_88));
	PE pe121_89(.x(x89),.w(w121_88),.acc(r121_88),.res(r121_89),.clk(clk),.wout(w121_89));
	PE pe121_90(.x(x90),.w(w121_89),.acc(r121_89),.res(r121_90),.clk(clk),.wout(w121_90));
	PE pe121_91(.x(x91),.w(w121_90),.acc(r121_90),.res(r121_91),.clk(clk),.wout(w121_91));
	PE pe121_92(.x(x92),.w(w121_91),.acc(r121_91),.res(r121_92),.clk(clk),.wout(w121_92));
	PE pe121_93(.x(x93),.w(w121_92),.acc(r121_92),.res(r121_93),.clk(clk),.wout(w121_93));
	PE pe121_94(.x(x94),.w(w121_93),.acc(r121_93),.res(r121_94),.clk(clk),.wout(w121_94));
	PE pe121_95(.x(x95),.w(w121_94),.acc(r121_94),.res(r121_95),.clk(clk),.wout(w121_95));
	PE pe121_96(.x(x96),.w(w121_95),.acc(r121_95),.res(r121_96),.clk(clk),.wout(w121_96));
	PE pe121_97(.x(x97),.w(w121_96),.acc(r121_96),.res(r121_97),.clk(clk),.wout(w121_97));
	PE pe121_98(.x(x98),.w(w121_97),.acc(r121_97),.res(r121_98),.clk(clk),.wout(w121_98));
	PE pe121_99(.x(x99),.w(w121_98),.acc(r121_98),.res(r121_99),.clk(clk),.wout(w121_99));
	PE pe121_100(.x(x100),.w(w121_99),.acc(r121_99),.res(r121_100),.clk(clk),.wout(w121_100));
	PE pe121_101(.x(x101),.w(w121_100),.acc(r121_100),.res(r121_101),.clk(clk),.wout(w121_101));
	PE pe121_102(.x(x102),.w(w121_101),.acc(r121_101),.res(r121_102),.clk(clk),.wout(w121_102));
	PE pe121_103(.x(x103),.w(w121_102),.acc(r121_102),.res(r121_103),.clk(clk),.wout(w121_103));
	PE pe121_104(.x(x104),.w(w121_103),.acc(r121_103),.res(r121_104),.clk(clk),.wout(w121_104));
	PE pe121_105(.x(x105),.w(w121_104),.acc(r121_104),.res(r121_105),.clk(clk),.wout(w121_105));
	PE pe121_106(.x(x106),.w(w121_105),.acc(r121_105),.res(r121_106),.clk(clk),.wout(w121_106));
	PE pe121_107(.x(x107),.w(w121_106),.acc(r121_106),.res(r121_107),.clk(clk),.wout(w121_107));
	PE pe121_108(.x(x108),.w(w121_107),.acc(r121_107),.res(r121_108),.clk(clk),.wout(w121_108));
	PE pe121_109(.x(x109),.w(w121_108),.acc(r121_108),.res(r121_109),.clk(clk),.wout(w121_109));
	PE pe121_110(.x(x110),.w(w121_109),.acc(r121_109),.res(r121_110),.clk(clk),.wout(w121_110));
	PE pe121_111(.x(x111),.w(w121_110),.acc(r121_110),.res(r121_111),.clk(clk),.wout(w121_111));
	PE pe121_112(.x(x112),.w(w121_111),.acc(r121_111),.res(r121_112),.clk(clk),.wout(w121_112));
	PE pe121_113(.x(x113),.w(w121_112),.acc(r121_112),.res(r121_113),.clk(clk),.wout(w121_113));
	PE pe121_114(.x(x114),.w(w121_113),.acc(r121_113),.res(r121_114),.clk(clk),.wout(w121_114));
	PE pe121_115(.x(x115),.w(w121_114),.acc(r121_114),.res(r121_115),.clk(clk),.wout(w121_115));
	PE pe121_116(.x(x116),.w(w121_115),.acc(r121_115),.res(r121_116),.clk(clk),.wout(w121_116));
	PE pe121_117(.x(x117),.w(w121_116),.acc(r121_116),.res(r121_117),.clk(clk),.wout(w121_117));
	PE pe121_118(.x(x118),.w(w121_117),.acc(r121_117),.res(r121_118),.clk(clk),.wout(w121_118));
	PE pe121_119(.x(x119),.w(w121_118),.acc(r121_118),.res(r121_119),.clk(clk),.wout(w121_119));
	PE pe121_120(.x(x120),.w(w121_119),.acc(r121_119),.res(r121_120),.clk(clk),.wout(w121_120));
	PE pe121_121(.x(x121),.w(w121_120),.acc(r121_120),.res(r121_121),.clk(clk),.wout(w121_121));
	PE pe121_122(.x(x122),.w(w121_121),.acc(r121_121),.res(r121_122),.clk(clk),.wout(w121_122));
	PE pe121_123(.x(x123),.w(w121_122),.acc(r121_122),.res(r121_123),.clk(clk),.wout(w121_123));
	PE pe121_124(.x(x124),.w(w121_123),.acc(r121_123),.res(r121_124),.clk(clk),.wout(w121_124));
	PE pe121_125(.x(x125),.w(w121_124),.acc(r121_124),.res(r121_125),.clk(clk),.wout(w121_125));
	PE pe121_126(.x(x126),.w(w121_125),.acc(r121_125),.res(r121_126),.clk(clk),.wout(w121_126));
	PE pe121_127(.x(x127),.w(w121_126),.acc(r121_126),.res(result121),.clk(clk),.wout(weight121));

	PE pe122_0(.x(x0),.w(w122),.acc(32'h0),.res(r122_0),.clk(clk),.wout(w122_0));
	PE pe122_1(.x(x1),.w(w122_0),.acc(r122_0),.res(r122_1),.clk(clk),.wout(w122_1));
	PE pe122_2(.x(x2),.w(w122_1),.acc(r122_1),.res(r122_2),.clk(clk),.wout(w122_2));
	PE pe122_3(.x(x3),.w(w122_2),.acc(r122_2),.res(r122_3),.clk(clk),.wout(w122_3));
	PE pe122_4(.x(x4),.w(w122_3),.acc(r122_3),.res(r122_4),.clk(clk),.wout(w122_4));
	PE pe122_5(.x(x5),.w(w122_4),.acc(r122_4),.res(r122_5),.clk(clk),.wout(w122_5));
	PE pe122_6(.x(x6),.w(w122_5),.acc(r122_5),.res(r122_6),.clk(clk),.wout(w122_6));
	PE pe122_7(.x(x7),.w(w122_6),.acc(r122_6),.res(r122_7),.clk(clk),.wout(w122_7));
	PE pe122_8(.x(x8),.w(w122_7),.acc(r122_7),.res(r122_8),.clk(clk),.wout(w122_8));
	PE pe122_9(.x(x9),.w(w122_8),.acc(r122_8),.res(r122_9),.clk(clk),.wout(w122_9));
	PE pe122_10(.x(x10),.w(w122_9),.acc(r122_9),.res(r122_10),.clk(clk),.wout(w122_10));
	PE pe122_11(.x(x11),.w(w122_10),.acc(r122_10),.res(r122_11),.clk(clk),.wout(w122_11));
	PE pe122_12(.x(x12),.w(w122_11),.acc(r122_11),.res(r122_12),.clk(clk),.wout(w122_12));
	PE pe122_13(.x(x13),.w(w122_12),.acc(r122_12),.res(r122_13),.clk(clk),.wout(w122_13));
	PE pe122_14(.x(x14),.w(w122_13),.acc(r122_13),.res(r122_14),.clk(clk),.wout(w122_14));
	PE pe122_15(.x(x15),.w(w122_14),.acc(r122_14),.res(r122_15),.clk(clk),.wout(w122_15));
	PE pe122_16(.x(x16),.w(w122_15),.acc(r122_15),.res(r122_16),.clk(clk),.wout(w122_16));
	PE pe122_17(.x(x17),.w(w122_16),.acc(r122_16),.res(r122_17),.clk(clk),.wout(w122_17));
	PE pe122_18(.x(x18),.w(w122_17),.acc(r122_17),.res(r122_18),.clk(clk),.wout(w122_18));
	PE pe122_19(.x(x19),.w(w122_18),.acc(r122_18),.res(r122_19),.clk(clk),.wout(w122_19));
	PE pe122_20(.x(x20),.w(w122_19),.acc(r122_19),.res(r122_20),.clk(clk),.wout(w122_20));
	PE pe122_21(.x(x21),.w(w122_20),.acc(r122_20),.res(r122_21),.clk(clk),.wout(w122_21));
	PE pe122_22(.x(x22),.w(w122_21),.acc(r122_21),.res(r122_22),.clk(clk),.wout(w122_22));
	PE pe122_23(.x(x23),.w(w122_22),.acc(r122_22),.res(r122_23),.clk(clk),.wout(w122_23));
	PE pe122_24(.x(x24),.w(w122_23),.acc(r122_23),.res(r122_24),.clk(clk),.wout(w122_24));
	PE pe122_25(.x(x25),.w(w122_24),.acc(r122_24),.res(r122_25),.clk(clk),.wout(w122_25));
	PE pe122_26(.x(x26),.w(w122_25),.acc(r122_25),.res(r122_26),.clk(clk),.wout(w122_26));
	PE pe122_27(.x(x27),.w(w122_26),.acc(r122_26),.res(r122_27),.clk(clk),.wout(w122_27));
	PE pe122_28(.x(x28),.w(w122_27),.acc(r122_27),.res(r122_28),.clk(clk),.wout(w122_28));
	PE pe122_29(.x(x29),.w(w122_28),.acc(r122_28),.res(r122_29),.clk(clk),.wout(w122_29));
	PE pe122_30(.x(x30),.w(w122_29),.acc(r122_29),.res(r122_30),.clk(clk),.wout(w122_30));
	PE pe122_31(.x(x31),.w(w122_30),.acc(r122_30),.res(r122_31),.clk(clk),.wout(w122_31));
	PE pe122_32(.x(x32),.w(w122_31),.acc(r122_31),.res(r122_32),.clk(clk),.wout(w122_32));
	PE pe122_33(.x(x33),.w(w122_32),.acc(r122_32),.res(r122_33),.clk(clk),.wout(w122_33));
	PE pe122_34(.x(x34),.w(w122_33),.acc(r122_33),.res(r122_34),.clk(clk),.wout(w122_34));
	PE pe122_35(.x(x35),.w(w122_34),.acc(r122_34),.res(r122_35),.clk(clk),.wout(w122_35));
	PE pe122_36(.x(x36),.w(w122_35),.acc(r122_35),.res(r122_36),.clk(clk),.wout(w122_36));
	PE pe122_37(.x(x37),.w(w122_36),.acc(r122_36),.res(r122_37),.clk(clk),.wout(w122_37));
	PE pe122_38(.x(x38),.w(w122_37),.acc(r122_37),.res(r122_38),.clk(clk),.wout(w122_38));
	PE pe122_39(.x(x39),.w(w122_38),.acc(r122_38),.res(r122_39),.clk(clk),.wout(w122_39));
	PE pe122_40(.x(x40),.w(w122_39),.acc(r122_39),.res(r122_40),.clk(clk),.wout(w122_40));
	PE pe122_41(.x(x41),.w(w122_40),.acc(r122_40),.res(r122_41),.clk(clk),.wout(w122_41));
	PE pe122_42(.x(x42),.w(w122_41),.acc(r122_41),.res(r122_42),.clk(clk),.wout(w122_42));
	PE pe122_43(.x(x43),.w(w122_42),.acc(r122_42),.res(r122_43),.clk(clk),.wout(w122_43));
	PE pe122_44(.x(x44),.w(w122_43),.acc(r122_43),.res(r122_44),.clk(clk),.wout(w122_44));
	PE pe122_45(.x(x45),.w(w122_44),.acc(r122_44),.res(r122_45),.clk(clk),.wout(w122_45));
	PE pe122_46(.x(x46),.w(w122_45),.acc(r122_45),.res(r122_46),.clk(clk),.wout(w122_46));
	PE pe122_47(.x(x47),.w(w122_46),.acc(r122_46),.res(r122_47),.clk(clk),.wout(w122_47));
	PE pe122_48(.x(x48),.w(w122_47),.acc(r122_47),.res(r122_48),.clk(clk),.wout(w122_48));
	PE pe122_49(.x(x49),.w(w122_48),.acc(r122_48),.res(r122_49),.clk(clk),.wout(w122_49));
	PE pe122_50(.x(x50),.w(w122_49),.acc(r122_49),.res(r122_50),.clk(clk),.wout(w122_50));
	PE pe122_51(.x(x51),.w(w122_50),.acc(r122_50),.res(r122_51),.clk(clk),.wout(w122_51));
	PE pe122_52(.x(x52),.w(w122_51),.acc(r122_51),.res(r122_52),.clk(clk),.wout(w122_52));
	PE pe122_53(.x(x53),.w(w122_52),.acc(r122_52),.res(r122_53),.clk(clk),.wout(w122_53));
	PE pe122_54(.x(x54),.w(w122_53),.acc(r122_53),.res(r122_54),.clk(clk),.wout(w122_54));
	PE pe122_55(.x(x55),.w(w122_54),.acc(r122_54),.res(r122_55),.clk(clk),.wout(w122_55));
	PE pe122_56(.x(x56),.w(w122_55),.acc(r122_55),.res(r122_56),.clk(clk),.wout(w122_56));
	PE pe122_57(.x(x57),.w(w122_56),.acc(r122_56),.res(r122_57),.clk(clk),.wout(w122_57));
	PE pe122_58(.x(x58),.w(w122_57),.acc(r122_57),.res(r122_58),.clk(clk),.wout(w122_58));
	PE pe122_59(.x(x59),.w(w122_58),.acc(r122_58),.res(r122_59),.clk(clk),.wout(w122_59));
	PE pe122_60(.x(x60),.w(w122_59),.acc(r122_59),.res(r122_60),.clk(clk),.wout(w122_60));
	PE pe122_61(.x(x61),.w(w122_60),.acc(r122_60),.res(r122_61),.clk(clk),.wout(w122_61));
	PE pe122_62(.x(x62),.w(w122_61),.acc(r122_61),.res(r122_62),.clk(clk),.wout(w122_62));
	PE pe122_63(.x(x63),.w(w122_62),.acc(r122_62),.res(r122_63),.clk(clk),.wout(w122_63));
	PE pe122_64(.x(x64),.w(w122_63),.acc(r122_63),.res(r122_64),.clk(clk),.wout(w122_64));
	PE pe122_65(.x(x65),.w(w122_64),.acc(r122_64),.res(r122_65),.clk(clk),.wout(w122_65));
	PE pe122_66(.x(x66),.w(w122_65),.acc(r122_65),.res(r122_66),.clk(clk),.wout(w122_66));
	PE pe122_67(.x(x67),.w(w122_66),.acc(r122_66),.res(r122_67),.clk(clk),.wout(w122_67));
	PE pe122_68(.x(x68),.w(w122_67),.acc(r122_67),.res(r122_68),.clk(clk),.wout(w122_68));
	PE pe122_69(.x(x69),.w(w122_68),.acc(r122_68),.res(r122_69),.clk(clk),.wout(w122_69));
	PE pe122_70(.x(x70),.w(w122_69),.acc(r122_69),.res(r122_70),.clk(clk),.wout(w122_70));
	PE pe122_71(.x(x71),.w(w122_70),.acc(r122_70),.res(r122_71),.clk(clk),.wout(w122_71));
	PE pe122_72(.x(x72),.w(w122_71),.acc(r122_71),.res(r122_72),.clk(clk),.wout(w122_72));
	PE pe122_73(.x(x73),.w(w122_72),.acc(r122_72),.res(r122_73),.clk(clk),.wout(w122_73));
	PE pe122_74(.x(x74),.w(w122_73),.acc(r122_73),.res(r122_74),.clk(clk),.wout(w122_74));
	PE pe122_75(.x(x75),.w(w122_74),.acc(r122_74),.res(r122_75),.clk(clk),.wout(w122_75));
	PE pe122_76(.x(x76),.w(w122_75),.acc(r122_75),.res(r122_76),.clk(clk),.wout(w122_76));
	PE pe122_77(.x(x77),.w(w122_76),.acc(r122_76),.res(r122_77),.clk(clk),.wout(w122_77));
	PE pe122_78(.x(x78),.w(w122_77),.acc(r122_77),.res(r122_78),.clk(clk),.wout(w122_78));
	PE pe122_79(.x(x79),.w(w122_78),.acc(r122_78),.res(r122_79),.clk(clk),.wout(w122_79));
	PE pe122_80(.x(x80),.w(w122_79),.acc(r122_79),.res(r122_80),.clk(clk),.wout(w122_80));
	PE pe122_81(.x(x81),.w(w122_80),.acc(r122_80),.res(r122_81),.clk(clk),.wout(w122_81));
	PE pe122_82(.x(x82),.w(w122_81),.acc(r122_81),.res(r122_82),.clk(clk),.wout(w122_82));
	PE pe122_83(.x(x83),.w(w122_82),.acc(r122_82),.res(r122_83),.clk(clk),.wout(w122_83));
	PE pe122_84(.x(x84),.w(w122_83),.acc(r122_83),.res(r122_84),.clk(clk),.wout(w122_84));
	PE pe122_85(.x(x85),.w(w122_84),.acc(r122_84),.res(r122_85),.clk(clk),.wout(w122_85));
	PE pe122_86(.x(x86),.w(w122_85),.acc(r122_85),.res(r122_86),.clk(clk),.wout(w122_86));
	PE pe122_87(.x(x87),.w(w122_86),.acc(r122_86),.res(r122_87),.clk(clk),.wout(w122_87));
	PE pe122_88(.x(x88),.w(w122_87),.acc(r122_87),.res(r122_88),.clk(clk),.wout(w122_88));
	PE pe122_89(.x(x89),.w(w122_88),.acc(r122_88),.res(r122_89),.clk(clk),.wout(w122_89));
	PE pe122_90(.x(x90),.w(w122_89),.acc(r122_89),.res(r122_90),.clk(clk),.wout(w122_90));
	PE pe122_91(.x(x91),.w(w122_90),.acc(r122_90),.res(r122_91),.clk(clk),.wout(w122_91));
	PE pe122_92(.x(x92),.w(w122_91),.acc(r122_91),.res(r122_92),.clk(clk),.wout(w122_92));
	PE pe122_93(.x(x93),.w(w122_92),.acc(r122_92),.res(r122_93),.clk(clk),.wout(w122_93));
	PE pe122_94(.x(x94),.w(w122_93),.acc(r122_93),.res(r122_94),.clk(clk),.wout(w122_94));
	PE pe122_95(.x(x95),.w(w122_94),.acc(r122_94),.res(r122_95),.clk(clk),.wout(w122_95));
	PE pe122_96(.x(x96),.w(w122_95),.acc(r122_95),.res(r122_96),.clk(clk),.wout(w122_96));
	PE pe122_97(.x(x97),.w(w122_96),.acc(r122_96),.res(r122_97),.clk(clk),.wout(w122_97));
	PE pe122_98(.x(x98),.w(w122_97),.acc(r122_97),.res(r122_98),.clk(clk),.wout(w122_98));
	PE pe122_99(.x(x99),.w(w122_98),.acc(r122_98),.res(r122_99),.clk(clk),.wout(w122_99));
	PE pe122_100(.x(x100),.w(w122_99),.acc(r122_99),.res(r122_100),.clk(clk),.wout(w122_100));
	PE pe122_101(.x(x101),.w(w122_100),.acc(r122_100),.res(r122_101),.clk(clk),.wout(w122_101));
	PE pe122_102(.x(x102),.w(w122_101),.acc(r122_101),.res(r122_102),.clk(clk),.wout(w122_102));
	PE pe122_103(.x(x103),.w(w122_102),.acc(r122_102),.res(r122_103),.clk(clk),.wout(w122_103));
	PE pe122_104(.x(x104),.w(w122_103),.acc(r122_103),.res(r122_104),.clk(clk),.wout(w122_104));
	PE pe122_105(.x(x105),.w(w122_104),.acc(r122_104),.res(r122_105),.clk(clk),.wout(w122_105));
	PE pe122_106(.x(x106),.w(w122_105),.acc(r122_105),.res(r122_106),.clk(clk),.wout(w122_106));
	PE pe122_107(.x(x107),.w(w122_106),.acc(r122_106),.res(r122_107),.clk(clk),.wout(w122_107));
	PE pe122_108(.x(x108),.w(w122_107),.acc(r122_107),.res(r122_108),.clk(clk),.wout(w122_108));
	PE pe122_109(.x(x109),.w(w122_108),.acc(r122_108),.res(r122_109),.clk(clk),.wout(w122_109));
	PE pe122_110(.x(x110),.w(w122_109),.acc(r122_109),.res(r122_110),.clk(clk),.wout(w122_110));
	PE pe122_111(.x(x111),.w(w122_110),.acc(r122_110),.res(r122_111),.clk(clk),.wout(w122_111));
	PE pe122_112(.x(x112),.w(w122_111),.acc(r122_111),.res(r122_112),.clk(clk),.wout(w122_112));
	PE pe122_113(.x(x113),.w(w122_112),.acc(r122_112),.res(r122_113),.clk(clk),.wout(w122_113));
	PE pe122_114(.x(x114),.w(w122_113),.acc(r122_113),.res(r122_114),.clk(clk),.wout(w122_114));
	PE pe122_115(.x(x115),.w(w122_114),.acc(r122_114),.res(r122_115),.clk(clk),.wout(w122_115));
	PE pe122_116(.x(x116),.w(w122_115),.acc(r122_115),.res(r122_116),.clk(clk),.wout(w122_116));
	PE pe122_117(.x(x117),.w(w122_116),.acc(r122_116),.res(r122_117),.clk(clk),.wout(w122_117));
	PE pe122_118(.x(x118),.w(w122_117),.acc(r122_117),.res(r122_118),.clk(clk),.wout(w122_118));
	PE pe122_119(.x(x119),.w(w122_118),.acc(r122_118),.res(r122_119),.clk(clk),.wout(w122_119));
	PE pe122_120(.x(x120),.w(w122_119),.acc(r122_119),.res(r122_120),.clk(clk),.wout(w122_120));
	PE pe122_121(.x(x121),.w(w122_120),.acc(r122_120),.res(r122_121),.clk(clk),.wout(w122_121));
	PE pe122_122(.x(x122),.w(w122_121),.acc(r122_121),.res(r122_122),.clk(clk),.wout(w122_122));
	PE pe122_123(.x(x123),.w(w122_122),.acc(r122_122),.res(r122_123),.clk(clk),.wout(w122_123));
	PE pe122_124(.x(x124),.w(w122_123),.acc(r122_123),.res(r122_124),.clk(clk),.wout(w122_124));
	PE pe122_125(.x(x125),.w(w122_124),.acc(r122_124),.res(r122_125),.clk(clk),.wout(w122_125));
	PE pe122_126(.x(x126),.w(w122_125),.acc(r122_125),.res(r122_126),.clk(clk),.wout(w122_126));
	PE pe122_127(.x(x127),.w(w122_126),.acc(r122_126),.res(result122),.clk(clk),.wout(weight122));

	PE pe123_0(.x(x0),.w(w123),.acc(32'h0),.res(r123_0),.clk(clk),.wout(w123_0));
	PE pe123_1(.x(x1),.w(w123_0),.acc(r123_0),.res(r123_1),.clk(clk),.wout(w123_1));
	PE pe123_2(.x(x2),.w(w123_1),.acc(r123_1),.res(r123_2),.clk(clk),.wout(w123_2));
	PE pe123_3(.x(x3),.w(w123_2),.acc(r123_2),.res(r123_3),.clk(clk),.wout(w123_3));
	PE pe123_4(.x(x4),.w(w123_3),.acc(r123_3),.res(r123_4),.clk(clk),.wout(w123_4));
	PE pe123_5(.x(x5),.w(w123_4),.acc(r123_4),.res(r123_5),.clk(clk),.wout(w123_5));
	PE pe123_6(.x(x6),.w(w123_5),.acc(r123_5),.res(r123_6),.clk(clk),.wout(w123_6));
	PE pe123_7(.x(x7),.w(w123_6),.acc(r123_6),.res(r123_7),.clk(clk),.wout(w123_7));
	PE pe123_8(.x(x8),.w(w123_7),.acc(r123_7),.res(r123_8),.clk(clk),.wout(w123_8));
	PE pe123_9(.x(x9),.w(w123_8),.acc(r123_8),.res(r123_9),.clk(clk),.wout(w123_9));
	PE pe123_10(.x(x10),.w(w123_9),.acc(r123_9),.res(r123_10),.clk(clk),.wout(w123_10));
	PE pe123_11(.x(x11),.w(w123_10),.acc(r123_10),.res(r123_11),.clk(clk),.wout(w123_11));
	PE pe123_12(.x(x12),.w(w123_11),.acc(r123_11),.res(r123_12),.clk(clk),.wout(w123_12));
	PE pe123_13(.x(x13),.w(w123_12),.acc(r123_12),.res(r123_13),.clk(clk),.wout(w123_13));
	PE pe123_14(.x(x14),.w(w123_13),.acc(r123_13),.res(r123_14),.clk(clk),.wout(w123_14));
	PE pe123_15(.x(x15),.w(w123_14),.acc(r123_14),.res(r123_15),.clk(clk),.wout(w123_15));
	PE pe123_16(.x(x16),.w(w123_15),.acc(r123_15),.res(r123_16),.clk(clk),.wout(w123_16));
	PE pe123_17(.x(x17),.w(w123_16),.acc(r123_16),.res(r123_17),.clk(clk),.wout(w123_17));
	PE pe123_18(.x(x18),.w(w123_17),.acc(r123_17),.res(r123_18),.clk(clk),.wout(w123_18));
	PE pe123_19(.x(x19),.w(w123_18),.acc(r123_18),.res(r123_19),.clk(clk),.wout(w123_19));
	PE pe123_20(.x(x20),.w(w123_19),.acc(r123_19),.res(r123_20),.clk(clk),.wout(w123_20));
	PE pe123_21(.x(x21),.w(w123_20),.acc(r123_20),.res(r123_21),.clk(clk),.wout(w123_21));
	PE pe123_22(.x(x22),.w(w123_21),.acc(r123_21),.res(r123_22),.clk(clk),.wout(w123_22));
	PE pe123_23(.x(x23),.w(w123_22),.acc(r123_22),.res(r123_23),.clk(clk),.wout(w123_23));
	PE pe123_24(.x(x24),.w(w123_23),.acc(r123_23),.res(r123_24),.clk(clk),.wout(w123_24));
	PE pe123_25(.x(x25),.w(w123_24),.acc(r123_24),.res(r123_25),.clk(clk),.wout(w123_25));
	PE pe123_26(.x(x26),.w(w123_25),.acc(r123_25),.res(r123_26),.clk(clk),.wout(w123_26));
	PE pe123_27(.x(x27),.w(w123_26),.acc(r123_26),.res(r123_27),.clk(clk),.wout(w123_27));
	PE pe123_28(.x(x28),.w(w123_27),.acc(r123_27),.res(r123_28),.clk(clk),.wout(w123_28));
	PE pe123_29(.x(x29),.w(w123_28),.acc(r123_28),.res(r123_29),.clk(clk),.wout(w123_29));
	PE pe123_30(.x(x30),.w(w123_29),.acc(r123_29),.res(r123_30),.clk(clk),.wout(w123_30));
	PE pe123_31(.x(x31),.w(w123_30),.acc(r123_30),.res(r123_31),.clk(clk),.wout(w123_31));
	PE pe123_32(.x(x32),.w(w123_31),.acc(r123_31),.res(r123_32),.clk(clk),.wout(w123_32));
	PE pe123_33(.x(x33),.w(w123_32),.acc(r123_32),.res(r123_33),.clk(clk),.wout(w123_33));
	PE pe123_34(.x(x34),.w(w123_33),.acc(r123_33),.res(r123_34),.clk(clk),.wout(w123_34));
	PE pe123_35(.x(x35),.w(w123_34),.acc(r123_34),.res(r123_35),.clk(clk),.wout(w123_35));
	PE pe123_36(.x(x36),.w(w123_35),.acc(r123_35),.res(r123_36),.clk(clk),.wout(w123_36));
	PE pe123_37(.x(x37),.w(w123_36),.acc(r123_36),.res(r123_37),.clk(clk),.wout(w123_37));
	PE pe123_38(.x(x38),.w(w123_37),.acc(r123_37),.res(r123_38),.clk(clk),.wout(w123_38));
	PE pe123_39(.x(x39),.w(w123_38),.acc(r123_38),.res(r123_39),.clk(clk),.wout(w123_39));
	PE pe123_40(.x(x40),.w(w123_39),.acc(r123_39),.res(r123_40),.clk(clk),.wout(w123_40));
	PE pe123_41(.x(x41),.w(w123_40),.acc(r123_40),.res(r123_41),.clk(clk),.wout(w123_41));
	PE pe123_42(.x(x42),.w(w123_41),.acc(r123_41),.res(r123_42),.clk(clk),.wout(w123_42));
	PE pe123_43(.x(x43),.w(w123_42),.acc(r123_42),.res(r123_43),.clk(clk),.wout(w123_43));
	PE pe123_44(.x(x44),.w(w123_43),.acc(r123_43),.res(r123_44),.clk(clk),.wout(w123_44));
	PE pe123_45(.x(x45),.w(w123_44),.acc(r123_44),.res(r123_45),.clk(clk),.wout(w123_45));
	PE pe123_46(.x(x46),.w(w123_45),.acc(r123_45),.res(r123_46),.clk(clk),.wout(w123_46));
	PE pe123_47(.x(x47),.w(w123_46),.acc(r123_46),.res(r123_47),.clk(clk),.wout(w123_47));
	PE pe123_48(.x(x48),.w(w123_47),.acc(r123_47),.res(r123_48),.clk(clk),.wout(w123_48));
	PE pe123_49(.x(x49),.w(w123_48),.acc(r123_48),.res(r123_49),.clk(clk),.wout(w123_49));
	PE pe123_50(.x(x50),.w(w123_49),.acc(r123_49),.res(r123_50),.clk(clk),.wout(w123_50));
	PE pe123_51(.x(x51),.w(w123_50),.acc(r123_50),.res(r123_51),.clk(clk),.wout(w123_51));
	PE pe123_52(.x(x52),.w(w123_51),.acc(r123_51),.res(r123_52),.clk(clk),.wout(w123_52));
	PE pe123_53(.x(x53),.w(w123_52),.acc(r123_52),.res(r123_53),.clk(clk),.wout(w123_53));
	PE pe123_54(.x(x54),.w(w123_53),.acc(r123_53),.res(r123_54),.clk(clk),.wout(w123_54));
	PE pe123_55(.x(x55),.w(w123_54),.acc(r123_54),.res(r123_55),.clk(clk),.wout(w123_55));
	PE pe123_56(.x(x56),.w(w123_55),.acc(r123_55),.res(r123_56),.clk(clk),.wout(w123_56));
	PE pe123_57(.x(x57),.w(w123_56),.acc(r123_56),.res(r123_57),.clk(clk),.wout(w123_57));
	PE pe123_58(.x(x58),.w(w123_57),.acc(r123_57),.res(r123_58),.clk(clk),.wout(w123_58));
	PE pe123_59(.x(x59),.w(w123_58),.acc(r123_58),.res(r123_59),.clk(clk),.wout(w123_59));
	PE pe123_60(.x(x60),.w(w123_59),.acc(r123_59),.res(r123_60),.clk(clk),.wout(w123_60));
	PE pe123_61(.x(x61),.w(w123_60),.acc(r123_60),.res(r123_61),.clk(clk),.wout(w123_61));
	PE pe123_62(.x(x62),.w(w123_61),.acc(r123_61),.res(r123_62),.clk(clk),.wout(w123_62));
	PE pe123_63(.x(x63),.w(w123_62),.acc(r123_62),.res(r123_63),.clk(clk),.wout(w123_63));
	PE pe123_64(.x(x64),.w(w123_63),.acc(r123_63),.res(r123_64),.clk(clk),.wout(w123_64));
	PE pe123_65(.x(x65),.w(w123_64),.acc(r123_64),.res(r123_65),.clk(clk),.wout(w123_65));
	PE pe123_66(.x(x66),.w(w123_65),.acc(r123_65),.res(r123_66),.clk(clk),.wout(w123_66));
	PE pe123_67(.x(x67),.w(w123_66),.acc(r123_66),.res(r123_67),.clk(clk),.wout(w123_67));
	PE pe123_68(.x(x68),.w(w123_67),.acc(r123_67),.res(r123_68),.clk(clk),.wout(w123_68));
	PE pe123_69(.x(x69),.w(w123_68),.acc(r123_68),.res(r123_69),.clk(clk),.wout(w123_69));
	PE pe123_70(.x(x70),.w(w123_69),.acc(r123_69),.res(r123_70),.clk(clk),.wout(w123_70));
	PE pe123_71(.x(x71),.w(w123_70),.acc(r123_70),.res(r123_71),.clk(clk),.wout(w123_71));
	PE pe123_72(.x(x72),.w(w123_71),.acc(r123_71),.res(r123_72),.clk(clk),.wout(w123_72));
	PE pe123_73(.x(x73),.w(w123_72),.acc(r123_72),.res(r123_73),.clk(clk),.wout(w123_73));
	PE pe123_74(.x(x74),.w(w123_73),.acc(r123_73),.res(r123_74),.clk(clk),.wout(w123_74));
	PE pe123_75(.x(x75),.w(w123_74),.acc(r123_74),.res(r123_75),.clk(clk),.wout(w123_75));
	PE pe123_76(.x(x76),.w(w123_75),.acc(r123_75),.res(r123_76),.clk(clk),.wout(w123_76));
	PE pe123_77(.x(x77),.w(w123_76),.acc(r123_76),.res(r123_77),.clk(clk),.wout(w123_77));
	PE pe123_78(.x(x78),.w(w123_77),.acc(r123_77),.res(r123_78),.clk(clk),.wout(w123_78));
	PE pe123_79(.x(x79),.w(w123_78),.acc(r123_78),.res(r123_79),.clk(clk),.wout(w123_79));
	PE pe123_80(.x(x80),.w(w123_79),.acc(r123_79),.res(r123_80),.clk(clk),.wout(w123_80));
	PE pe123_81(.x(x81),.w(w123_80),.acc(r123_80),.res(r123_81),.clk(clk),.wout(w123_81));
	PE pe123_82(.x(x82),.w(w123_81),.acc(r123_81),.res(r123_82),.clk(clk),.wout(w123_82));
	PE pe123_83(.x(x83),.w(w123_82),.acc(r123_82),.res(r123_83),.clk(clk),.wout(w123_83));
	PE pe123_84(.x(x84),.w(w123_83),.acc(r123_83),.res(r123_84),.clk(clk),.wout(w123_84));
	PE pe123_85(.x(x85),.w(w123_84),.acc(r123_84),.res(r123_85),.clk(clk),.wout(w123_85));
	PE pe123_86(.x(x86),.w(w123_85),.acc(r123_85),.res(r123_86),.clk(clk),.wout(w123_86));
	PE pe123_87(.x(x87),.w(w123_86),.acc(r123_86),.res(r123_87),.clk(clk),.wout(w123_87));
	PE pe123_88(.x(x88),.w(w123_87),.acc(r123_87),.res(r123_88),.clk(clk),.wout(w123_88));
	PE pe123_89(.x(x89),.w(w123_88),.acc(r123_88),.res(r123_89),.clk(clk),.wout(w123_89));
	PE pe123_90(.x(x90),.w(w123_89),.acc(r123_89),.res(r123_90),.clk(clk),.wout(w123_90));
	PE pe123_91(.x(x91),.w(w123_90),.acc(r123_90),.res(r123_91),.clk(clk),.wout(w123_91));
	PE pe123_92(.x(x92),.w(w123_91),.acc(r123_91),.res(r123_92),.clk(clk),.wout(w123_92));
	PE pe123_93(.x(x93),.w(w123_92),.acc(r123_92),.res(r123_93),.clk(clk),.wout(w123_93));
	PE pe123_94(.x(x94),.w(w123_93),.acc(r123_93),.res(r123_94),.clk(clk),.wout(w123_94));
	PE pe123_95(.x(x95),.w(w123_94),.acc(r123_94),.res(r123_95),.clk(clk),.wout(w123_95));
	PE pe123_96(.x(x96),.w(w123_95),.acc(r123_95),.res(r123_96),.clk(clk),.wout(w123_96));
	PE pe123_97(.x(x97),.w(w123_96),.acc(r123_96),.res(r123_97),.clk(clk),.wout(w123_97));
	PE pe123_98(.x(x98),.w(w123_97),.acc(r123_97),.res(r123_98),.clk(clk),.wout(w123_98));
	PE pe123_99(.x(x99),.w(w123_98),.acc(r123_98),.res(r123_99),.clk(clk),.wout(w123_99));
	PE pe123_100(.x(x100),.w(w123_99),.acc(r123_99),.res(r123_100),.clk(clk),.wout(w123_100));
	PE pe123_101(.x(x101),.w(w123_100),.acc(r123_100),.res(r123_101),.clk(clk),.wout(w123_101));
	PE pe123_102(.x(x102),.w(w123_101),.acc(r123_101),.res(r123_102),.clk(clk),.wout(w123_102));
	PE pe123_103(.x(x103),.w(w123_102),.acc(r123_102),.res(r123_103),.clk(clk),.wout(w123_103));
	PE pe123_104(.x(x104),.w(w123_103),.acc(r123_103),.res(r123_104),.clk(clk),.wout(w123_104));
	PE pe123_105(.x(x105),.w(w123_104),.acc(r123_104),.res(r123_105),.clk(clk),.wout(w123_105));
	PE pe123_106(.x(x106),.w(w123_105),.acc(r123_105),.res(r123_106),.clk(clk),.wout(w123_106));
	PE pe123_107(.x(x107),.w(w123_106),.acc(r123_106),.res(r123_107),.clk(clk),.wout(w123_107));
	PE pe123_108(.x(x108),.w(w123_107),.acc(r123_107),.res(r123_108),.clk(clk),.wout(w123_108));
	PE pe123_109(.x(x109),.w(w123_108),.acc(r123_108),.res(r123_109),.clk(clk),.wout(w123_109));
	PE pe123_110(.x(x110),.w(w123_109),.acc(r123_109),.res(r123_110),.clk(clk),.wout(w123_110));
	PE pe123_111(.x(x111),.w(w123_110),.acc(r123_110),.res(r123_111),.clk(clk),.wout(w123_111));
	PE pe123_112(.x(x112),.w(w123_111),.acc(r123_111),.res(r123_112),.clk(clk),.wout(w123_112));
	PE pe123_113(.x(x113),.w(w123_112),.acc(r123_112),.res(r123_113),.clk(clk),.wout(w123_113));
	PE pe123_114(.x(x114),.w(w123_113),.acc(r123_113),.res(r123_114),.clk(clk),.wout(w123_114));
	PE pe123_115(.x(x115),.w(w123_114),.acc(r123_114),.res(r123_115),.clk(clk),.wout(w123_115));
	PE pe123_116(.x(x116),.w(w123_115),.acc(r123_115),.res(r123_116),.clk(clk),.wout(w123_116));
	PE pe123_117(.x(x117),.w(w123_116),.acc(r123_116),.res(r123_117),.clk(clk),.wout(w123_117));
	PE pe123_118(.x(x118),.w(w123_117),.acc(r123_117),.res(r123_118),.clk(clk),.wout(w123_118));
	PE pe123_119(.x(x119),.w(w123_118),.acc(r123_118),.res(r123_119),.clk(clk),.wout(w123_119));
	PE pe123_120(.x(x120),.w(w123_119),.acc(r123_119),.res(r123_120),.clk(clk),.wout(w123_120));
	PE pe123_121(.x(x121),.w(w123_120),.acc(r123_120),.res(r123_121),.clk(clk),.wout(w123_121));
	PE pe123_122(.x(x122),.w(w123_121),.acc(r123_121),.res(r123_122),.clk(clk),.wout(w123_122));
	PE pe123_123(.x(x123),.w(w123_122),.acc(r123_122),.res(r123_123),.clk(clk),.wout(w123_123));
	PE pe123_124(.x(x124),.w(w123_123),.acc(r123_123),.res(r123_124),.clk(clk),.wout(w123_124));
	PE pe123_125(.x(x125),.w(w123_124),.acc(r123_124),.res(r123_125),.clk(clk),.wout(w123_125));
	PE pe123_126(.x(x126),.w(w123_125),.acc(r123_125),.res(r123_126),.clk(clk),.wout(w123_126));
	PE pe123_127(.x(x127),.w(w123_126),.acc(r123_126),.res(result123),.clk(clk),.wout(weight123));

	PE pe124_0(.x(x0),.w(w124),.acc(32'h0),.res(r124_0),.clk(clk),.wout(w124_0));
	PE pe124_1(.x(x1),.w(w124_0),.acc(r124_0),.res(r124_1),.clk(clk),.wout(w124_1));
	PE pe124_2(.x(x2),.w(w124_1),.acc(r124_1),.res(r124_2),.clk(clk),.wout(w124_2));
	PE pe124_3(.x(x3),.w(w124_2),.acc(r124_2),.res(r124_3),.clk(clk),.wout(w124_3));
	PE pe124_4(.x(x4),.w(w124_3),.acc(r124_3),.res(r124_4),.clk(clk),.wout(w124_4));
	PE pe124_5(.x(x5),.w(w124_4),.acc(r124_4),.res(r124_5),.clk(clk),.wout(w124_5));
	PE pe124_6(.x(x6),.w(w124_5),.acc(r124_5),.res(r124_6),.clk(clk),.wout(w124_6));
	PE pe124_7(.x(x7),.w(w124_6),.acc(r124_6),.res(r124_7),.clk(clk),.wout(w124_7));
	PE pe124_8(.x(x8),.w(w124_7),.acc(r124_7),.res(r124_8),.clk(clk),.wout(w124_8));
	PE pe124_9(.x(x9),.w(w124_8),.acc(r124_8),.res(r124_9),.clk(clk),.wout(w124_9));
	PE pe124_10(.x(x10),.w(w124_9),.acc(r124_9),.res(r124_10),.clk(clk),.wout(w124_10));
	PE pe124_11(.x(x11),.w(w124_10),.acc(r124_10),.res(r124_11),.clk(clk),.wout(w124_11));
	PE pe124_12(.x(x12),.w(w124_11),.acc(r124_11),.res(r124_12),.clk(clk),.wout(w124_12));
	PE pe124_13(.x(x13),.w(w124_12),.acc(r124_12),.res(r124_13),.clk(clk),.wout(w124_13));
	PE pe124_14(.x(x14),.w(w124_13),.acc(r124_13),.res(r124_14),.clk(clk),.wout(w124_14));
	PE pe124_15(.x(x15),.w(w124_14),.acc(r124_14),.res(r124_15),.clk(clk),.wout(w124_15));
	PE pe124_16(.x(x16),.w(w124_15),.acc(r124_15),.res(r124_16),.clk(clk),.wout(w124_16));
	PE pe124_17(.x(x17),.w(w124_16),.acc(r124_16),.res(r124_17),.clk(clk),.wout(w124_17));
	PE pe124_18(.x(x18),.w(w124_17),.acc(r124_17),.res(r124_18),.clk(clk),.wout(w124_18));
	PE pe124_19(.x(x19),.w(w124_18),.acc(r124_18),.res(r124_19),.clk(clk),.wout(w124_19));
	PE pe124_20(.x(x20),.w(w124_19),.acc(r124_19),.res(r124_20),.clk(clk),.wout(w124_20));
	PE pe124_21(.x(x21),.w(w124_20),.acc(r124_20),.res(r124_21),.clk(clk),.wout(w124_21));
	PE pe124_22(.x(x22),.w(w124_21),.acc(r124_21),.res(r124_22),.clk(clk),.wout(w124_22));
	PE pe124_23(.x(x23),.w(w124_22),.acc(r124_22),.res(r124_23),.clk(clk),.wout(w124_23));
	PE pe124_24(.x(x24),.w(w124_23),.acc(r124_23),.res(r124_24),.clk(clk),.wout(w124_24));
	PE pe124_25(.x(x25),.w(w124_24),.acc(r124_24),.res(r124_25),.clk(clk),.wout(w124_25));
	PE pe124_26(.x(x26),.w(w124_25),.acc(r124_25),.res(r124_26),.clk(clk),.wout(w124_26));
	PE pe124_27(.x(x27),.w(w124_26),.acc(r124_26),.res(r124_27),.clk(clk),.wout(w124_27));
	PE pe124_28(.x(x28),.w(w124_27),.acc(r124_27),.res(r124_28),.clk(clk),.wout(w124_28));
	PE pe124_29(.x(x29),.w(w124_28),.acc(r124_28),.res(r124_29),.clk(clk),.wout(w124_29));
	PE pe124_30(.x(x30),.w(w124_29),.acc(r124_29),.res(r124_30),.clk(clk),.wout(w124_30));
	PE pe124_31(.x(x31),.w(w124_30),.acc(r124_30),.res(r124_31),.clk(clk),.wout(w124_31));
	PE pe124_32(.x(x32),.w(w124_31),.acc(r124_31),.res(r124_32),.clk(clk),.wout(w124_32));
	PE pe124_33(.x(x33),.w(w124_32),.acc(r124_32),.res(r124_33),.clk(clk),.wout(w124_33));
	PE pe124_34(.x(x34),.w(w124_33),.acc(r124_33),.res(r124_34),.clk(clk),.wout(w124_34));
	PE pe124_35(.x(x35),.w(w124_34),.acc(r124_34),.res(r124_35),.clk(clk),.wout(w124_35));
	PE pe124_36(.x(x36),.w(w124_35),.acc(r124_35),.res(r124_36),.clk(clk),.wout(w124_36));
	PE pe124_37(.x(x37),.w(w124_36),.acc(r124_36),.res(r124_37),.clk(clk),.wout(w124_37));
	PE pe124_38(.x(x38),.w(w124_37),.acc(r124_37),.res(r124_38),.clk(clk),.wout(w124_38));
	PE pe124_39(.x(x39),.w(w124_38),.acc(r124_38),.res(r124_39),.clk(clk),.wout(w124_39));
	PE pe124_40(.x(x40),.w(w124_39),.acc(r124_39),.res(r124_40),.clk(clk),.wout(w124_40));
	PE pe124_41(.x(x41),.w(w124_40),.acc(r124_40),.res(r124_41),.clk(clk),.wout(w124_41));
	PE pe124_42(.x(x42),.w(w124_41),.acc(r124_41),.res(r124_42),.clk(clk),.wout(w124_42));
	PE pe124_43(.x(x43),.w(w124_42),.acc(r124_42),.res(r124_43),.clk(clk),.wout(w124_43));
	PE pe124_44(.x(x44),.w(w124_43),.acc(r124_43),.res(r124_44),.clk(clk),.wout(w124_44));
	PE pe124_45(.x(x45),.w(w124_44),.acc(r124_44),.res(r124_45),.clk(clk),.wout(w124_45));
	PE pe124_46(.x(x46),.w(w124_45),.acc(r124_45),.res(r124_46),.clk(clk),.wout(w124_46));
	PE pe124_47(.x(x47),.w(w124_46),.acc(r124_46),.res(r124_47),.clk(clk),.wout(w124_47));
	PE pe124_48(.x(x48),.w(w124_47),.acc(r124_47),.res(r124_48),.clk(clk),.wout(w124_48));
	PE pe124_49(.x(x49),.w(w124_48),.acc(r124_48),.res(r124_49),.clk(clk),.wout(w124_49));
	PE pe124_50(.x(x50),.w(w124_49),.acc(r124_49),.res(r124_50),.clk(clk),.wout(w124_50));
	PE pe124_51(.x(x51),.w(w124_50),.acc(r124_50),.res(r124_51),.clk(clk),.wout(w124_51));
	PE pe124_52(.x(x52),.w(w124_51),.acc(r124_51),.res(r124_52),.clk(clk),.wout(w124_52));
	PE pe124_53(.x(x53),.w(w124_52),.acc(r124_52),.res(r124_53),.clk(clk),.wout(w124_53));
	PE pe124_54(.x(x54),.w(w124_53),.acc(r124_53),.res(r124_54),.clk(clk),.wout(w124_54));
	PE pe124_55(.x(x55),.w(w124_54),.acc(r124_54),.res(r124_55),.clk(clk),.wout(w124_55));
	PE pe124_56(.x(x56),.w(w124_55),.acc(r124_55),.res(r124_56),.clk(clk),.wout(w124_56));
	PE pe124_57(.x(x57),.w(w124_56),.acc(r124_56),.res(r124_57),.clk(clk),.wout(w124_57));
	PE pe124_58(.x(x58),.w(w124_57),.acc(r124_57),.res(r124_58),.clk(clk),.wout(w124_58));
	PE pe124_59(.x(x59),.w(w124_58),.acc(r124_58),.res(r124_59),.clk(clk),.wout(w124_59));
	PE pe124_60(.x(x60),.w(w124_59),.acc(r124_59),.res(r124_60),.clk(clk),.wout(w124_60));
	PE pe124_61(.x(x61),.w(w124_60),.acc(r124_60),.res(r124_61),.clk(clk),.wout(w124_61));
	PE pe124_62(.x(x62),.w(w124_61),.acc(r124_61),.res(r124_62),.clk(clk),.wout(w124_62));
	PE pe124_63(.x(x63),.w(w124_62),.acc(r124_62),.res(r124_63),.clk(clk),.wout(w124_63));
	PE pe124_64(.x(x64),.w(w124_63),.acc(r124_63),.res(r124_64),.clk(clk),.wout(w124_64));
	PE pe124_65(.x(x65),.w(w124_64),.acc(r124_64),.res(r124_65),.clk(clk),.wout(w124_65));
	PE pe124_66(.x(x66),.w(w124_65),.acc(r124_65),.res(r124_66),.clk(clk),.wout(w124_66));
	PE pe124_67(.x(x67),.w(w124_66),.acc(r124_66),.res(r124_67),.clk(clk),.wout(w124_67));
	PE pe124_68(.x(x68),.w(w124_67),.acc(r124_67),.res(r124_68),.clk(clk),.wout(w124_68));
	PE pe124_69(.x(x69),.w(w124_68),.acc(r124_68),.res(r124_69),.clk(clk),.wout(w124_69));
	PE pe124_70(.x(x70),.w(w124_69),.acc(r124_69),.res(r124_70),.clk(clk),.wout(w124_70));
	PE pe124_71(.x(x71),.w(w124_70),.acc(r124_70),.res(r124_71),.clk(clk),.wout(w124_71));
	PE pe124_72(.x(x72),.w(w124_71),.acc(r124_71),.res(r124_72),.clk(clk),.wout(w124_72));
	PE pe124_73(.x(x73),.w(w124_72),.acc(r124_72),.res(r124_73),.clk(clk),.wout(w124_73));
	PE pe124_74(.x(x74),.w(w124_73),.acc(r124_73),.res(r124_74),.clk(clk),.wout(w124_74));
	PE pe124_75(.x(x75),.w(w124_74),.acc(r124_74),.res(r124_75),.clk(clk),.wout(w124_75));
	PE pe124_76(.x(x76),.w(w124_75),.acc(r124_75),.res(r124_76),.clk(clk),.wout(w124_76));
	PE pe124_77(.x(x77),.w(w124_76),.acc(r124_76),.res(r124_77),.clk(clk),.wout(w124_77));
	PE pe124_78(.x(x78),.w(w124_77),.acc(r124_77),.res(r124_78),.clk(clk),.wout(w124_78));
	PE pe124_79(.x(x79),.w(w124_78),.acc(r124_78),.res(r124_79),.clk(clk),.wout(w124_79));
	PE pe124_80(.x(x80),.w(w124_79),.acc(r124_79),.res(r124_80),.clk(clk),.wout(w124_80));
	PE pe124_81(.x(x81),.w(w124_80),.acc(r124_80),.res(r124_81),.clk(clk),.wout(w124_81));
	PE pe124_82(.x(x82),.w(w124_81),.acc(r124_81),.res(r124_82),.clk(clk),.wout(w124_82));
	PE pe124_83(.x(x83),.w(w124_82),.acc(r124_82),.res(r124_83),.clk(clk),.wout(w124_83));
	PE pe124_84(.x(x84),.w(w124_83),.acc(r124_83),.res(r124_84),.clk(clk),.wout(w124_84));
	PE pe124_85(.x(x85),.w(w124_84),.acc(r124_84),.res(r124_85),.clk(clk),.wout(w124_85));
	PE pe124_86(.x(x86),.w(w124_85),.acc(r124_85),.res(r124_86),.clk(clk),.wout(w124_86));
	PE pe124_87(.x(x87),.w(w124_86),.acc(r124_86),.res(r124_87),.clk(clk),.wout(w124_87));
	PE pe124_88(.x(x88),.w(w124_87),.acc(r124_87),.res(r124_88),.clk(clk),.wout(w124_88));
	PE pe124_89(.x(x89),.w(w124_88),.acc(r124_88),.res(r124_89),.clk(clk),.wout(w124_89));
	PE pe124_90(.x(x90),.w(w124_89),.acc(r124_89),.res(r124_90),.clk(clk),.wout(w124_90));
	PE pe124_91(.x(x91),.w(w124_90),.acc(r124_90),.res(r124_91),.clk(clk),.wout(w124_91));
	PE pe124_92(.x(x92),.w(w124_91),.acc(r124_91),.res(r124_92),.clk(clk),.wout(w124_92));
	PE pe124_93(.x(x93),.w(w124_92),.acc(r124_92),.res(r124_93),.clk(clk),.wout(w124_93));
	PE pe124_94(.x(x94),.w(w124_93),.acc(r124_93),.res(r124_94),.clk(clk),.wout(w124_94));
	PE pe124_95(.x(x95),.w(w124_94),.acc(r124_94),.res(r124_95),.clk(clk),.wout(w124_95));
	PE pe124_96(.x(x96),.w(w124_95),.acc(r124_95),.res(r124_96),.clk(clk),.wout(w124_96));
	PE pe124_97(.x(x97),.w(w124_96),.acc(r124_96),.res(r124_97),.clk(clk),.wout(w124_97));
	PE pe124_98(.x(x98),.w(w124_97),.acc(r124_97),.res(r124_98),.clk(clk),.wout(w124_98));
	PE pe124_99(.x(x99),.w(w124_98),.acc(r124_98),.res(r124_99),.clk(clk),.wout(w124_99));
	PE pe124_100(.x(x100),.w(w124_99),.acc(r124_99),.res(r124_100),.clk(clk),.wout(w124_100));
	PE pe124_101(.x(x101),.w(w124_100),.acc(r124_100),.res(r124_101),.clk(clk),.wout(w124_101));
	PE pe124_102(.x(x102),.w(w124_101),.acc(r124_101),.res(r124_102),.clk(clk),.wout(w124_102));
	PE pe124_103(.x(x103),.w(w124_102),.acc(r124_102),.res(r124_103),.clk(clk),.wout(w124_103));
	PE pe124_104(.x(x104),.w(w124_103),.acc(r124_103),.res(r124_104),.clk(clk),.wout(w124_104));
	PE pe124_105(.x(x105),.w(w124_104),.acc(r124_104),.res(r124_105),.clk(clk),.wout(w124_105));
	PE pe124_106(.x(x106),.w(w124_105),.acc(r124_105),.res(r124_106),.clk(clk),.wout(w124_106));
	PE pe124_107(.x(x107),.w(w124_106),.acc(r124_106),.res(r124_107),.clk(clk),.wout(w124_107));
	PE pe124_108(.x(x108),.w(w124_107),.acc(r124_107),.res(r124_108),.clk(clk),.wout(w124_108));
	PE pe124_109(.x(x109),.w(w124_108),.acc(r124_108),.res(r124_109),.clk(clk),.wout(w124_109));
	PE pe124_110(.x(x110),.w(w124_109),.acc(r124_109),.res(r124_110),.clk(clk),.wout(w124_110));
	PE pe124_111(.x(x111),.w(w124_110),.acc(r124_110),.res(r124_111),.clk(clk),.wout(w124_111));
	PE pe124_112(.x(x112),.w(w124_111),.acc(r124_111),.res(r124_112),.clk(clk),.wout(w124_112));
	PE pe124_113(.x(x113),.w(w124_112),.acc(r124_112),.res(r124_113),.clk(clk),.wout(w124_113));
	PE pe124_114(.x(x114),.w(w124_113),.acc(r124_113),.res(r124_114),.clk(clk),.wout(w124_114));
	PE pe124_115(.x(x115),.w(w124_114),.acc(r124_114),.res(r124_115),.clk(clk),.wout(w124_115));
	PE pe124_116(.x(x116),.w(w124_115),.acc(r124_115),.res(r124_116),.clk(clk),.wout(w124_116));
	PE pe124_117(.x(x117),.w(w124_116),.acc(r124_116),.res(r124_117),.clk(clk),.wout(w124_117));
	PE pe124_118(.x(x118),.w(w124_117),.acc(r124_117),.res(r124_118),.clk(clk),.wout(w124_118));
	PE pe124_119(.x(x119),.w(w124_118),.acc(r124_118),.res(r124_119),.clk(clk),.wout(w124_119));
	PE pe124_120(.x(x120),.w(w124_119),.acc(r124_119),.res(r124_120),.clk(clk),.wout(w124_120));
	PE pe124_121(.x(x121),.w(w124_120),.acc(r124_120),.res(r124_121),.clk(clk),.wout(w124_121));
	PE pe124_122(.x(x122),.w(w124_121),.acc(r124_121),.res(r124_122),.clk(clk),.wout(w124_122));
	PE pe124_123(.x(x123),.w(w124_122),.acc(r124_122),.res(r124_123),.clk(clk),.wout(w124_123));
	PE pe124_124(.x(x124),.w(w124_123),.acc(r124_123),.res(r124_124),.clk(clk),.wout(w124_124));
	PE pe124_125(.x(x125),.w(w124_124),.acc(r124_124),.res(r124_125),.clk(clk),.wout(w124_125));
	PE pe124_126(.x(x126),.w(w124_125),.acc(r124_125),.res(r124_126),.clk(clk),.wout(w124_126));
	PE pe124_127(.x(x127),.w(w124_126),.acc(r124_126),.res(result124),.clk(clk),.wout(weight124));

	PE pe125_0(.x(x0),.w(w125),.acc(32'h0),.res(r125_0),.clk(clk),.wout(w125_0));
	PE pe125_1(.x(x1),.w(w125_0),.acc(r125_0),.res(r125_1),.clk(clk),.wout(w125_1));
	PE pe125_2(.x(x2),.w(w125_1),.acc(r125_1),.res(r125_2),.clk(clk),.wout(w125_2));
	PE pe125_3(.x(x3),.w(w125_2),.acc(r125_2),.res(r125_3),.clk(clk),.wout(w125_3));
	PE pe125_4(.x(x4),.w(w125_3),.acc(r125_3),.res(r125_4),.clk(clk),.wout(w125_4));
	PE pe125_5(.x(x5),.w(w125_4),.acc(r125_4),.res(r125_5),.clk(clk),.wout(w125_5));
	PE pe125_6(.x(x6),.w(w125_5),.acc(r125_5),.res(r125_6),.clk(clk),.wout(w125_6));
	PE pe125_7(.x(x7),.w(w125_6),.acc(r125_6),.res(r125_7),.clk(clk),.wout(w125_7));
	PE pe125_8(.x(x8),.w(w125_7),.acc(r125_7),.res(r125_8),.clk(clk),.wout(w125_8));
	PE pe125_9(.x(x9),.w(w125_8),.acc(r125_8),.res(r125_9),.clk(clk),.wout(w125_9));
	PE pe125_10(.x(x10),.w(w125_9),.acc(r125_9),.res(r125_10),.clk(clk),.wout(w125_10));
	PE pe125_11(.x(x11),.w(w125_10),.acc(r125_10),.res(r125_11),.clk(clk),.wout(w125_11));
	PE pe125_12(.x(x12),.w(w125_11),.acc(r125_11),.res(r125_12),.clk(clk),.wout(w125_12));
	PE pe125_13(.x(x13),.w(w125_12),.acc(r125_12),.res(r125_13),.clk(clk),.wout(w125_13));
	PE pe125_14(.x(x14),.w(w125_13),.acc(r125_13),.res(r125_14),.clk(clk),.wout(w125_14));
	PE pe125_15(.x(x15),.w(w125_14),.acc(r125_14),.res(r125_15),.clk(clk),.wout(w125_15));
	PE pe125_16(.x(x16),.w(w125_15),.acc(r125_15),.res(r125_16),.clk(clk),.wout(w125_16));
	PE pe125_17(.x(x17),.w(w125_16),.acc(r125_16),.res(r125_17),.clk(clk),.wout(w125_17));
	PE pe125_18(.x(x18),.w(w125_17),.acc(r125_17),.res(r125_18),.clk(clk),.wout(w125_18));
	PE pe125_19(.x(x19),.w(w125_18),.acc(r125_18),.res(r125_19),.clk(clk),.wout(w125_19));
	PE pe125_20(.x(x20),.w(w125_19),.acc(r125_19),.res(r125_20),.clk(clk),.wout(w125_20));
	PE pe125_21(.x(x21),.w(w125_20),.acc(r125_20),.res(r125_21),.clk(clk),.wout(w125_21));
	PE pe125_22(.x(x22),.w(w125_21),.acc(r125_21),.res(r125_22),.clk(clk),.wout(w125_22));
	PE pe125_23(.x(x23),.w(w125_22),.acc(r125_22),.res(r125_23),.clk(clk),.wout(w125_23));
	PE pe125_24(.x(x24),.w(w125_23),.acc(r125_23),.res(r125_24),.clk(clk),.wout(w125_24));
	PE pe125_25(.x(x25),.w(w125_24),.acc(r125_24),.res(r125_25),.clk(clk),.wout(w125_25));
	PE pe125_26(.x(x26),.w(w125_25),.acc(r125_25),.res(r125_26),.clk(clk),.wout(w125_26));
	PE pe125_27(.x(x27),.w(w125_26),.acc(r125_26),.res(r125_27),.clk(clk),.wout(w125_27));
	PE pe125_28(.x(x28),.w(w125_27),.acc(r125_27),.res(r125_28),.clk(clk),.wout(w125_28));
	PE pe125_29(.x(x29),.w(w125_28),.acc(r125_28),.res(r125_29),.clk(clk),.wout(w125_29));
	PE pe125_30(.x(x30),.w(w125_29),.acc(r125_29),.res(r125_30),.clk(clk),.wout(w125_30));
	PE pe125_31(.x(x31),.w(w125_30),.acc(r125_30),.res(r125_31),.clk(clk),.wout(w125_31));
	PE pe125_32(.x(x32),.w(w125_31),.acc(r125_31),.res(r125_32),.clk(clk),.wout(w125_32));
	PE pe125_33(.x(x33),.w(w125_32),.acc(r125_32),.res(r125_33),.clk(clk),.wout(w125_33));
	PE pe125_34(.x(x34),.w(w125_33),.acc(r125_33),.res(r125_34),.clk(clk),.wout(w125_34));
	PE pe125_35(.x(x35),.w(w125_34),.acc(r125_34),.res(r125_35),.clk(clk),.wout(w125_35));
	PE pe125_36(.x(x36),.w(w125_35),.acc(r125_35),.res(r125_36),.clk(clk),.wout(w125_36));
	PE pe125_37(.x(x37),.w(w125_36),.acc(r125_36),.res(r125_37),.clk(clk),.wout(w125_37));
	PE pe125_38(.x(x38),.w(w125_37),.acc(r125_37),.res(r125_38),.clk(clk),.wout(w125_38));
	PE pe125_39(.x(x39),.w(w125_38),.acc(r125_38),.res(r125_39),.clk(clk),.wout(w125_39));
	PE pe125_40(.x(x40),.w(w125_39),.acc(r125_39),.res(r125_40),.clk(clk),.wout(w125_40));
	PE pe125_41(.x(x41),.w(w125_40),.acc(r125_40),.res(r125_41),.clk(clk),.wout(w125_41));
	PE pe125_42(.x(x42),.w(w125_41),.acc(r125_41),.res(r125_42),.clk(clk),.wout(w125_42));
	PE pe125_43(.x(x43),.w(w125_42),.acc(r125_42),.res(r125_43),.clk(clk),.wout(w125_43));
	PE pe125_44(.x(x44),.w(w125_43),.acc(r125_43),.res(r125_44),.clk(clk),.wout(w125_44));
	PE pe125_45(.x(x45),.w(w125_44),.acc(r125_44),.res(r125_45),.clk(clk),.wout(w125_45));
	PE pe125_46(.x(x46),.w(w125_45),.acc(r125_45),.res(r125_46),.clk(clk),.wout(w125_46));
	PE pe125_47(.x(x47),.w(w125_46),.acc(r125_46),.res(r125_47),.clk(clk),.wout(w125_47));
	PE pe125_48(.x(x48),.w(w125_47),.acc(r125_47),.res(r125_48),.clk(clk),.wout(w125_48));
	PE pe125_49(.x(x49),.w(w125_48),.acc(r125_48),.res(r125_49),.clk(clk),.wout(w125_49));
	PE pe125_50(.x(x50),.w(w125_49),.acc(r125_49),.res(r125_50),.clk(clk),.wout(w125_50));
	PE pe125_51(.x(x51),.w(w125_50),.acc(r125_50),.res(r125_51),.clk(clk),.wout(w125_51));
	PE pe125_52(.x(x52),.w(w125_51),.acc(r125_51),.res(r125_52),.clk(clk),.wout(w125_52));
	PE pe125_53(.x(x53),.w(w125_52),.acc(r125_52),.res(r125_53),.clk(clk),.wout(w125_53));
	PE pe125_54(.x(x54),.w(w125_53),.acc(r125_53),.res(r125_54),.clk(clk),.wout(w125_54));
	PE pe125_55(.x(x55),.w(w125_54),.acc(r125_54),.res(r125_55),.clk(clk),.wout(w125_55));
	PE pe125_56(.x(x56),.w(w125_55),.acc(r125_55),.res(r125_56),.clk(clk),.wout(w125_56));
	PE pe125_57(.x(x57),.w(w125_56),.acc(r125_56),.res(r125_57),.clk(clk),.wout(w125_57));
	PE pe125_58(.x(x58),.w(w125_57),.acc(r125_57),.res(r125_58),.clk(clk),.wout(w125_58));
	PE pe125_59(.x(x59),.w(w125_58),.acc(r125_58),.res(r125_59),.clk(clk),.wout(w125_59));
	PE pe125_60(.x(x60),.w(w125_59),.acc(r125_59),.res(r125_60),.clk(clk),.wout(w125_60));
	PE pe125_61(.x(x61),.w(w125_60),.acc(r125_60),.res(r125_61),.clk(clk),.wout(w125_61));
	PE pe125_62(.x(x62),.w(w125_61),.acc(r125_61),.res(r125_62),.clk(clk),.wout(w125_62));
	PE pe125_63(.x(x63),.w(w125_62),.acc(r125_62),.res(r125_63),.clk(clk),.wout(w125_63));
	PE pe125_64(.x(x64),.w(w125_63),.acc(r125_63),.res(r125_64),.clk(clk),.wout(w125_64));
	PE pe125_65(.x(x65),.w(w125_64),.acc(r125_64),.res(r125_65),.clk(clk),.wout(w125_65));
	PE pe125_66(.x(x66),.w(w125_65),.acc(r125_65),.res(r125_66),.clk(clk),.wout(w125_66));
	PE pe125_67(.x(x67),.w(w125_66),.acc(r125_66),.res(r125_67),.clk(clk),.wout(w125_67));
	PE pe125_68(.x(x68),.w(w125_67),.acc(r125_67),.res(r125_68),.clk(clk),.wout(w125_68));
	PE pe125_69(.x(x69),.w(w125_68),.acc(r125_68),.res(r125_69),.clk(clk),.wout(w125_69));
	PE pe125_70(.x(x70),.w(w125_69),.acc(r125_69),.res(r125_70),.clk(clk),.wout(w125_70));
	PE pe125_71(.x(x71),.w(w125_70),.acc(r125_70),.res(r125_71),.clk(clk),.wout(w125_71));
	PE pe125_72(.x(x72),.w(w125_71),.acc(r125_71),.res(r125_72),.clk(clk),.wout(w125_72));
	PE pe125_73(.x(x73),.w(w125_72),.acc(r125_72),.res(r125_73),.clk(clk),.wout(w125_73));
	PE pe125_74(.x(x74),.w(w125_73),.acc(r125_73),.res(r125_74),.clk(clk),.wout(w125_74));
	PE pe125_75(.x(x75),.w(w125_74),.acc(r125_74),.res(r125_75),.clk(clk),.wout(w125_75));
	PE pe125_76(.x(x76),.w(w125_75),.acc(r125_75),.res(r125_76),.clk(clk),.wout(w125_76));
	PE pe125_77(.x(x77),.w(w125_76),.acc(r125_76),.res(r125_77),.clk(clk),.wout(w125_77));
	PE pe125_78(.x(x78),.w(w125_77),.acc(r125_77),.res(r125_78),.clk(clk),.wout(w125_78));
	PE pe125_79(.x(x79),.w(w125_78),.acc(r125_78),.res(r125_79),.clk(clk),.wout(w125_79));
	PE pe125_80(.x(x80),.w(w125_79),.acc(r125_79),.res(r125_80),.clk(clk),.wout(w125_80));
	PE pe125_81(.x(x81),.w(w125_80),.acc(r125_80),.res(r125_81),.clk(clk),.wout(w125_81));
	PE pe125_82(.x(x82),.w(w125_81),.acc(r125_81),.res(r125_82),.clk(clk),.wout(w125_82));
	PE pe125_83(.x(x83),.w(w125_82),.acc(r125_82),.res(r125_83),.clk(clk),.wout(w125_83));
	PE pe125_84(.x(x84),.w(w125_83),.acc(r125_83),.res(r125_84),.clk(clk),.wout(w125_84));
	PE pe125_85(.x(x85),.w(w125_84),.acc(r125_84),.res(r125_85),.clk(clk),.wout(w125_85));
	PE pe125_86(.x(x86),.w(w125_85),.acc(r125_85),.res(r125_86),.clk(clk),.wout(w125_86));
	PE pe125_87(.x(x87),.w(w125_86),.acc(r125_86),.res(r125_87),.clk(clk),.wout(w125_87));
	PE pe125_88(.x(x88),.w(w125_87),.acc(r125_87),.res(r125_88),.clk(clk),.wout(w125_88));
	PE pe125_89(.x(x89),.w(w125_88),.acc(r125_88),.res(r125_89),.clk(clk),.wout(w125_89));
	PE pe125_90(.x(x90),.w(w125_89),.acc(r125_89),.res(r125_90),.clk(clk),.wout(w125_90));
	PE pe125_91(.x(x91),.w(w125_90),.acc(r125_90),.res(r125_91),.clk(clk),.wout(w125_91));
	PE pe125_92(.x(x92),.w(w125_91),.acc(r125_91),.res(r125_92),.clk(clk),.wout(w125_92));
	PE pe125_93(.x(x93),.w(w125_92),.acc(r125_92),.res(r125_93),.clk(clk),.wout(w125_93));
	PE pe125_94(.x(x94),.w(w125_93),.acc(r125_93),.res(r125_94),.clk(clk),.wout(w125_94));
	PE pe125_95(.x(x95),.w(w125_94),.acc(r125_94),.res(r125_95),.clk(clk),.wout(w125_95));
	PE pe125_96(.x(x96),.w(w125_95),.acc(r125_95),.res(r125_96),.clk(clk),.wout(w125_96));
	PE pe125_97(.x(x97),.w(w125_96),.acc(r125_96),.res(r125_97),.clk(clk),.wout(w125_97));
	PE pe125_98(.x(x98),.w(w125_97),.acc(r125_97),.res(r125_98),.clk(clk),.wout(w125_98));
	PE pe125_99(.x(x99),.w(w125_98),.acc(r125_98),.res(r125_99),.clk(clk),.wout(w125_99));
	PE pe125_100(.x(x100),.w(w125_99),.acc(r125_99),.res(r125_100),.clk(clk),.wout(w125_100));
	PE pe125_101(.x(x101),.w(w125_100),.acc(r125_100),.res(r125_101),.clk(clk),.wout(w125_101));
	PE pe125_102(.x(x102),.w(w125_101),.acc(r125_101),.res(r125_102),.clk(clk),.wout(w125_102));
	PE pe125_103(.x(x103),.w(w125_102),.acc(r125_102),.res(r125_103),.clk(clk),.wout(w125_103));
	PE pe125_104(.x(x104),.w(w125_103),.acc(r125_103),.res(r125_104),.clk(clk),.wout(w125_104));
	PE pe125_105(.x(x105),.w(w125_104),.acc(r125_104),.res(r125_105),.clk(clk),.wout(w125_105));
	PE pe125_106(.x(x106),.w(w125_105),.acc(r125_105),.res(r125_106),.clk(clk),.wout(w125_106));
	PE pe125_107(.x(x107),.w(w125_106),.acc(r125_106),.res(r125_107),.clk(clk),.wout(w125_107));
	PE pe125_108(.x(x108),.w(w125_107),.acc(r125_107),.res(r125_108),.clk(clk),.wout(w125_108));
	PE pe125_109(.x(x109),.w(w125_108),.acc(r125_108),.res(r125_109),.clk(clk),.wout(w125_109));
	PE pe125_110(.x(x110),.w(w125_109),.acc(r125_109),.res(r125_110),.clk(clk),.wout(w125_110));
	PE pe125_111(.x(x111),.w(w125_110),.acc(r125_110),.res(r125_111),.clk(clk),.wout(w125_111));
	PE pe125_112(.x(x112),.w(w125_111),.acc(r125_111),.res(r125_112),.clk(clk),.wout(w125_112));
	PE pe125_113(.x(x113),.w(w125_112),.acc(r125_112),.res(r125_113),.clk(clk),.wout(w125_113));
	PE pe125_114(.x(x114),.w(w125_113),.acc(r125_113),.res(r125_114),.clk(clk),.wout(w125_114));
	PE pe125_115(.x(x115),.w(w125_114),.acc(r125_114),.res(r125_115),.clk(clk),.wout(w125_115));
	PE pe125_116(.x(x116),.w(w125_115),.acc(r125_115),.res(r125_116),.clk(clk),.wout(w125_116));
	PE pe125_117(.x(x117),.w(w125_116),.acc(r125_116),.res(r125_117),.clk(clk),.wout(w125_117));
	PE pe125_118(.x(x118),.w(w125_117),.acc(r125_117),.res(r125_118),.clk(clk),.wout(w125_118));
	PE pe125_119(.x(x119),.w(w125_118),.acc(r125_118),.res(r125_119),.clk(clk),.wout(w125_119));
	PE pe125_120(.x(x120),.w(w125_119),.acc(r125_119),.res(r125_120),.clk(clk),.wout(w125_120));
	PE pe125_121(.x(x121),.w(w125_120),.acc(r125_120),.res(r125_121),.clk(clk),.wout(w125_121));
	PE pe125_122(.x(x122),.w(w125_121),.acc(r125_121),.res(r125_122),.clk(clk),.wout(w125_122));
	PE pe125_123(.x(x123),.w(w125_122),.acc(r125_122),.res(r125_123),.clk(clk),.wout(w125_123));
	PE pe125_124(.x(x124),.w(w125_123),.acc(r125_123),.res(r125_124),.clk(clk),.wout(w125_124));
	PE pe125_125(.x(x125),.w(w125_124),.acc(r125_124),.res(r125_125),.clk(clk),.wout(w125_125));
	PE pe125_126(.x(x126),.w(w125_125),.acc(r125_125),.res(r125_126),.clk(clk),.wout(w125_126));
	PE pe125_127(.x(x127),.w(w125_126),.acc(r125_126),.res(result125),.clk(clk),.wout(weight125));

	PE pe126_0(.x(x0),.w(w126),.acc(32'h0),.res(r126_0),.clk(clk),.wout(w126_0));
	PE pe126_1(.x(x1),.w(w126_0),.acc(r126_0),.res(r126_1),.clk(clk),.wout(w126_1));
	PE pe126_2(.x(x2),.w(w126_1),.acc(r126_1),.res(r126_2),.clk(clk),.wout(w126_2));
	PE pe126_3(.x(x3),.w(w126_2),.acc(r126_2),.res(r126_3),.clk(clk),.wout(w126_3));
	PE pe126_4(.x(x4),.w(w126_3),.acc(r126_3),.res(r126_4),.clk(clk),.wout(w126_4));
	PE pe126_5(.x(x5),.w(w126_4),.acc(r126_4),.res(r126_5),.clk(clk),.wout(w126_5));
	PE pe126_6(.x(x6),.w(w126_5),.acc(r126_5),.res(r126_6),.clk(clk),.wout(w126_6));
	PE pe126_7(.x(x7),.w(w126_6),.acc(r126_6),.res(r126_7),.clk(clk),.wout(w126_7));
	PE pe126_8(.x(x8),.w(w126_7),.acc(r126_7),.res(r126_8),.clk(clk),.wout(w126_8));
	PE pe126_9(.x(x9),.w(w126_8),.acc(r126_8),.res(r126_9),.clk(clk),.wout(w126_9));
	PE pe126_10(.x(x10),.w(w126_9),.acc(r126_9),.res(r126_10),.clk(clk),.wout(w126_10));
	PE pe126_11(.x(x11),.w(w126_10),.acc(r126_10),.res(r126_11),.clk(clk),.wout(w126_11));
	PE pe126_12(.x(x12),.w(w126_11),.acc(r126_11),.res(r126_12),.clk(clk),.wout(w126_12));
	PE pe126_13(.x(x13),.w(w126_12),.acc(r126_12),.res(r126_13),.clk(clk),.wout(w126_13));
	PE pe126_14(.x(x14),.w(w126_13),.acc(r126_13),.res(r126_14),.clk(clk),.wout(w126_14));
	PE pe126_15(.x(x15),.w(w126_14),.acc(r126_14),.res(r126_15),.clk(clk),.wout(w126_15));
	PE pe126_16(.x(x16),.w(w126_15),.acc(r126_15),.res(r126_16),.clk(clk),.wout(w126_16));
	PE pe126_17(.x(x17),.w(w126_16),.acc(r126_16),.res(r126_17),.clk(clk),.wout(w126_17));
	PE pe126_18(.x(x18),.w(w126_17),.acc(r126_17),.res(r126_18),.clk(clk),.wout(w126_18));
	PE pe126_19(.x(x19),.w(w126_18),.acc(r126_18),.res(r126_19),.clk(clk),.wout(w126_19));
	PE pe126_20(.x(x20),.w(w126_19),.acc(r126_19),.res(r126_20),.clk(clk),.wout(w126_20));
	PE pe126_21(.x(x21),.w(w126_20),.acc(r126_20),.res(r126_21),.clk(clk),.wout(w126_21));
	PE pe126_22(.x(x22),.w(w126_21),.acc(r126_21),.res(r126_22),.clk(clk),.wout(w126_22));
	PE pe126_23(.x(x23),.w(w126_22),.acc(r126_22),.res(r126_23),.clk(clk),.wout(w126_23));
	PE pe126_24(.x(x24),.w(w126_23),.acc(r126_23),.res(r126_24),.clk(clk),.wout(w126_24));
	PE pe126_25(.x(x25),.w(w126_24),.acc(r126_24),.res(r126_25),.clk(clk),.wout(w126_25));
	PE pe126_26(.x(x26),.w(w126_25),.acc(r126_25),.res(r126_26),.clk(clk),.wout(w126_26));
	PE pe126_27(.x(x27),.w(w126_26),.acc(r126_26),.res(r126_27),.clk(clk),.wout(w126_27));
	PE pe126_28(.x(x28),.w(w126_27),.acc(r126_27),.res(r126_28),.clk(clk),.wout(w126_28));
	PE pe126_29(.x(x29),.w(w126_28),.acc(r126_28),.res(r126_29),.clk(clk),.wout(w126_29));
	PE pe126_30(.x(x30),.w(w126_29),.acc(r126_29),.res(r126_30),.clk(clk),.wout(w126_30));
	PE pe126_31(.x(x31),.w(w126_30),.acc(r126_30),.res(r126_31),.clk(clk),.wout(w126_31));
	PE pe126_32(.x(x32),.w(w126_31),.acc(r126_31),.res(r126_32),.clk(clk),.wout(w126_32));
	PE pe126_33(.x(x33),.w(w126_32),.acc(r126_32),.res(r126_33),.clk(clk),.wout(w126_33));
	PE pe126_34(.x(x34),.w(w126_33),.acc(r126_33),.res(r126_34),.clk(clk),.wout(w126_34));
	PE pe126_35(.x(x35),.w(w126_34),.acc(r126_34),.res(r126_35),.clk(clk),.wout(w126_35));
	PE pe126_36(.x(x36),.w(w126_35),.acc(r126_35),.res(r126_36),.clk(clk),.wout(w126_36));
	PE pe126_37(.x(x37),.w(w126_36),.acc(r126_36),.res(r126_37),.clk(clk),.wout(w126_37));
	PE pe126_38(.x(x38),.w(w126_37),.acc(r126_37),.res(r126_38),.clk(clk),.wout(w126_38));
	PE pe126_39(.x(x39),.w(w126_38),.acc(r126_38),.res(r126_39),.clk(clk),.wout(w126_39));
	PE pe126_40(.x(x40),.w(w126_39),.acc(r126_39),.res(r126_40),.clk(clk),.wout(w126_40));
	PE pe126_41(.x(x41),.w(w126_40),.acc(r126_40),.res(r126_41),.clk(clk),.wout(w126_41));
	PE pe126_42(.x(x42),.w(w126_41),.acc(r126_41),.res(r126_42),.clk(clk),.wout(w126_42));
	PE pe126_43(.x(x43),.w(w126_42),.acc(r126_42),.res(r126_43),.clk(clk),.wout(w126_43));
	PE pe126_44(.x(x44),.w(w126_43),.acc(r126_43),.res(r126_44),.clk(clk),.wout(w126_44));
	PE pe126_45(.x(x45),.w(w126_44),.acc(r126_44),.res(r126_45),.clk(clk),.wout(w126_45));
	PE pe126_46(.x(x46),.w(w126_45),.acc(r126_45),.res(r126_46),.clk(clk),.wout(w126_46));
	PE pe126_47(.x(x47),.w(w126_46),.acc(r126_46),.res(r126_47),.clk(clk),.wout(w126_47));
	PE pe126_48(.x(x48),.w(w126_47),.acc(r126_47),.res(r126_48),.clk(clk),.wout(w126_48));
	PE pe126_49(.x(x49),.w(w126_48),.acc(r126_48),.res(r126_49),.clk(clk),.wout(w126_49));
	PE pe126_50(.x(x50),.w(w126_49),.acc(r126_49),.res(r126_50),.clk(clk),.wout(w126_50));
	PE pe126_51(.x(x51),.w(w126_50),.acc(r126_50),.res(r126_51),.clk(clk),.wout(w126_51));
	PE pe126_52(.x(x52),.w(w126_51),.acc(r126_51),.res(r126_52),.clk(clk),.wout(w126_52));
	PE pe126_53(.x(x53),.w(w126_52),.acc(r126_52),.res(r126_53),.clk(clk),.wout(w126_53));
	PE pe126_54(.x(x54),.w(w126_53),.acc(r126_53),.res(r126_54),.clk(clk),.wout(w126_54));
	PE pe126_55(.x(x55),.w(w126_54),.acc(r126_54),.res(r126_55),.clk(clk),.wout(w126_55));
	PE pe126_56(.x(x56),.w(w126_55),.acc(r126_55),.res(r126_56),.clk(clk),.wout(w126_56));
	PE pe126_57(.x(x57),.w(w126_56),.acc(r126_56),.res(r126_57),.clk(clk),.wout(w126_57));
	PE pe126_58(.x(x58),.w(w126_57),.acc(r126_57),.res(r126_58),.clk(clk),.wout(w126_58));
	PE pe126_59(.x(x59),.w(w126_58),.acc(r126_58),.res(r126_59),.clk(clk),.wout(w126_59));
	PE pe126_60(.x(x60),.w(w126_59),.acc(r126_59),.res(r126_60),.clk(clk),.wout(w126_60));
	PE pe126_61(.x(x61),.w(w126_60),.acc(r126_60),.res(r126_61),.clk(clk),.wout(w126_61));
	PE pe126_62(.x(x62),.w(w126_61),.acc(r126_61),.res(r126_62),.clk(clk),.wout(w126_62));
	PE pe126_63(.x(x63),.w(w126_62),.acc(r126_62),.res(r126_63),.clk(clk),.wout(w126_63));
	PE pe126_64(.x(x64),.w(w126_63),.acc(r126_63),.res(r126_64),.clk(clk),.wout(w126_64));
	PE pe126_65(.x(x65),.w(w126_64),.acc(r126_64),.res(r126_65),.clk(clk),.wout(w126_65));
	PE pe126_66(.x(x66),.w(w126_65),.acc(r126_65),.res(r126_66),.clk(clk),.wout(w126_66));
	PE pe126_67(.x(x67),.w(w126_66),.acc(r126_66),.res(r126_67),.clk(clk),.wout(w126_67));
	PE pe126_68(.x(x68),.w(w126_67),.acc(r126_67),.res(r126_68),.clk(clk),.wout(w126_68));
	PE pe126_69(.x(x69),.w(w126_68),.acc(r126_68),.res(r126_69),.clk(clk),.wout(w126_69));
	PE pe126_70(.x(x70),.w(w126_69),.acc(r126_69),.res(r126_70),.clk(clk),.wout(w126_70));
	PE pe126_71(.x(x71),.w(w126_70),.acc(r126_70),.res(r126_71),.clk(clk),.wout(w126_71));
	PE pe126_72(.x(x72),.w(w126_71),.acc(r126_71),.res(r126_72),.clk(clk),.wout(w126_72));
	PE pe126_73(.x(x73),.w(w126_72),.acc(r126_72),.res(r126_73),.clk(clk),.wout(w126_73));
	PE pe126_74(.x(x74),.w(w126_73),.acc(r126_73),.res(r126_74),.clk(clk),.wout(w126_74));
	PE pe126_75(.x(x75),.w(w126_74),.acc(r126_74),.res(r126_75),.clk(clk),.wout(w126_75));
	PE pe126_76(.x(x76),.w(w126_75),.acc(r126_75),.res(r126_76),.clk(clk),.wout(w126_76));
	PE pe126_77(.x(x77),.w(w126_76),.acc(r126_76),.res(r126_77),.clk(clk),.wout(w126_77));
	PE pe126_78(.x(x78),.w(w126_77),.acc(r126_77),.res(r126_78),.clk(clk),.wout(w126_78));
	PE pe126_79(.x(x79),.w(w126_78),.acc(r126_78),.res(r126_79),.clk(clk),.wout(w126_79));
	PE pe126_80(.x(x80),.w(w126_79),.acc(r126_79),.res(r126_80),.clk(clk),.wout(w126_80));
	PE pe126_81(.x(x81),.w(w126_80),.acc(r126_80),.res(r126_81),.clk(clk),.wout(w126_81));
	PE pe126_82(.x(x82),.w(w126_81),.acc(r126_81),.res(r126_82),.clk(clk),.wout(w126_82));
	PE pe126_83(.x(x83),.w(w126_82),.acc(r126_82),.res(r126_83),.clk(clk),.wout(w126_83));
	PE pe126_84(.x(x84),.w(w126_83),.acc(r126_83),.res(r126_84),.clk(clk),.wout(w126_84));
	PE pe126_85(.x(x85),.w(w126_84),.acc(r126_84),.res(r126_85),.clk(clk),.wout(w126_85));
	PE pe126_86(.x(x86),.w(w126_85),.acc(r126_85),.res(r126_86),.clk(clk),.wout(w126_86));
	PE pe126_87(.x(x87),.w(w126_86),.acc(r126_86),.res(r126_87),.clk(clk),.wout(w126_87));
	PE pe126_88(.x(x88),.w(w126_87),.acc(r126_87),.res(r126_88),.clk(clk),.wout(w126_88));
	PE pe126_89(.x(x89),.w(w126_88),.acc(r126_88),.res(r126_89),.clk(clk),.wout(w126_89));
	PE pe126_90(.x(x90),.w(w126_89),.acc(r126_89),.res(r126_90),.clk(clk),.wout(w126_90));
	PE pe126_91(.x(x91),.w(w126_90),.acc(r126_90),.res(r126_91),.clk(clk),.wout(w126_91));
	PE pe126_92(.x(x92),.w(w126_91),.acc(r126_91),.res(r126_92),.clk(clk),.wout(w126_92));
	PE pe126_93(.x(x93),.w(w126_92),.acc(r126_92),.res(r126_93),.clk(clk),.wout(w126_93));
	PE pe126_94(.x(x94),.w(w126_93),.acc(r126_93),.res(r126_94),.clk(clk),.wout(w126_94));
	PE pe126_95(.x(x95),.w(w126_94),.acc(r126_94),.res(r126_95),.clk(clk),.wout(w126_95));
	PE pe126_96(.x(x96),.w(w126_95),.acc(r126_95),.res(r126_96),.clk(clk),.wout(w126_96));
	PE pe126_97(.x(x97),.w(w126_96),.acc(r126_96),.res(r126_97),.clk(clk),.wout(w126_97));
	PE pe126_98(.x(x98),.w(w126_97),.acc(r126_97),.res(r126_98),.clk(clk),.wout(w126_98));
	PE pe126_99(.x(x99),.w(w126_98),.acc(r126_98),.res(r126_99),.clk(clk),.wout(w126_99));
	PE pe126_100(.x(x100),.w(w126_99),.acc(r126_99),.res(r126_100),.clk(clk),.wout(w126_100));
	PE pe126_101(.x(x101),.w(w126_100),.acc(r126_100),.res(r126_101),.clk(clk),.wout(w126_101));
	PE pe126_102(.x(x102),.w(w126_101),.acc(r126_101),.res(r126_102),.clk(clk),.wout(w126_102));
	PE pe126_103(.x(x103),.w(w126_102),.acc(r126_102),.res(r126_103),.clk(clk),.wout(w126_103));
	PE pe126_104(.x(x104),.w(w126_103),.acc(r126_103),.res(r126_104),.clk(clk),.wout(w126_104));
	PE pe126_105(.x(x105),.w(w126_104),.acc(r126_104),.res(r126_105),.clk(clk),.wout(w126_105));
	PE pe126_106(.x(x106),.w(w126_105),.acc(r126_105),.res(r126_106),.clk(clk),.wout(w126_106));
	PE pe126_107(.x(x107),.w(w126_106),.acc(r126_106),.res(r126_107),.clk(clk),.wout(w126_107));
	PE pe126_108(.x(x108),.w(w126_107),.acc(r126_107),.res(r126_108),.clk(clk),.wout(w126_108));
	PE pe126_109(.x(x109),.w(w126_108),.acc(r126_108),.res(r126_109),.clk(clk),.wout(w126_109));
	PE pe126_110(.x(x110),.w(w126_109),.acc(r126_109),.res(r126_110),.clk(clk),.wout(w126_110));
	PE pe126_111(.x(x111),.w(w126_110),.acc(r126_110),.res(r126_111),.clk(clk),.wout(w126_111));
	PE pe126_112(.x(x112),.w(w126_111),.acc(r126_111),.res(r126_112),.clk(clk),.wout(w126_112));
	PE pe126_113(.x(x113),.w(w126_112),.acc(r126_112),.res(r126_113),.clk(clk),.wout(w126_113));
	PE pe126_114(.x(x114),.w(w126_113),.acc(r126_113),.res(r126_114),.clk(clk),.wout(w126_114));
	PE pe126_115(.x(x115),.w(w126_114),.acc(r126_114),.res(r126_115),.clk(clk),.wout(w126_115));
	PE pe126_116(.x(x116),.w(w126_115),.acc(r126_115),.res(r126_116),.clk(clk),.wout(w126_116));
	PE pe126_117(.x(x117),.w(w126_116),.acc(r126_116),.res(r126_117),.clk(clk),.wout(w126_117));
	PE pe126_118(.x(x118),.w(w126_117),.acc(r126_117),.res(r126_118),.clk(clk),.wout(w126_118));
	PE pe126_119(.x(x119),.w(w126_118),.acc(r126_118),.res(r126_119),.clk(clk),.wout(w126_119));
	PE pe126_120(.x(x120),.w(w126_119),.acc(r126_119),.res(r126_120),.clk(clk),.wout(w126_120));
	PE pe126_121(.x(x121),.w(w126_120),.acc(r126_120),.res(r126_121),.clk(clk),.wout(w126_121));
	PE pe126_122(.x(x122),.w(w126_121),.acc(r126_121),.res(r126_122),.clk(clk),.wout(w126_122));
	PE pe126_123(.x(x123),.w(w126_122),.acc(r126_122),.res(r126_123),.clk(clk),.wout(w126_123));
	PE pe126_124(.x(x124),.w(w126_123),.acc(r126_123),.res(r126_124),.clk(clk),.wout(w126_124));
	PE pe126_125(.x(x125),.w(w126_124),.acc(r126_124),.res(r126_125),.clk(clk),.wout(w126_125));
	PE pe126_126(.x(x126),.w(w126_125),.acc(r126_125),.res(r126_126),.clk(clk),.wout(w126_126));
	PE pe126_127(.x(x127),.w(w126_126),.acc(r126_126),.res(result126),.clk(clk),.wout(weight126));

	PE_syn pe127_0(.x(x0),.w(w127),.acc(32'h0),.res(r127_0),.clk(clk),.wout(w127_0));
	PE pe127_1(.x(x1),.w(w127_0),.acc(r127_0),.res(r127_1),.clk(clk),.wout(w127_1));
	PE pe127_2(.x(x2),.w(w127_1),.acc(r127_1),.res(r127_2),.clk(clk),.wout(w127_2));
	PE pe127_3(.x(x3),.w(w127_2),.acc(r127_2),.res(r127_3),.clk(clk),.wout(w127_3));
	PE pe127_4(.x(x4),.w(w127_3),.acc(r127_3),.res(r127_4),.clk(clk),.wout(w127_4));
	PE pe127_5(.x(x5),.w(w127_4),.acc(r127_4),.res(r127_5),.clk(clk),.wout(w127_5));
	PE pe127_6(.x(x6),.w(w127_5),.acc(r127_5),.res(r127_6),.clk(clk),.wout(w127_6));
	PE pe127_7(.x(x7),.w(w127_6),.acc(r127_6),.res(r127_7),.clk(clk),.wout(w127_7));
	PE pe127_8(.x(x8),.w(w127_7),.acc(r127_7),.res(r127_8),.clk(clk),.wout(w127_8));
	PE pe127_9(.x(x9),.w(w127_8),.acc(r127_8),.res(r127_9),.clk(clk),.wout(w127_9));
	PE pe127_10(.x(x10),.w(w127_9),.acc(r127_9),.res(r127_10),.clk(clk),.wout(w127_10));
	PE pe127_11(.x(x11),.w(w127_10),.acc(r127_10),.res(r127_11),.clk(clk),.wout(w127_11));
	PE pe127_12(.x(x12),.w(w127_11),.acc(r127_11),.res(r127_12),.clk(clk),.wout(w127_12));
	PE pe127_13(.x(x13),.w(w127_12),.acc(r127_12),.res(r127_13),.clk(clk),.wout(w127_13));
	PE pe127_14(.x(x14),.w(w127_13),.acc(r127_13),.res(r127_14),.clk(clk),.wout(w127_14));
	PE pe127_15(.x(x15),.w(w127_14),.acc(r127_14),.res(r127_15),.clk(clk),.wout(w127_15));
	PE pe127_16(.x(x16),.w(w127_15),.acc(r127_15),.res(r127_16),.clk(clk),.wout(w127_16));
	PE pe127_17(.x(x17),.w(w127_16),.acc(r127_16),.res(r127_17),.clk(clk),.wout(w127_17));
	PE pe127_18(.x(x18),.w(w127_17),.acc(r127_17),.res(r127_18),.clk(clk),.wout(w127_18));
	PE pe127_19(.x(x19),.w(w127_18),.acc(r127_18),.res(r127_19),.clk(clk),.wout(w127_19));
	PE pe127_20(.x(x20),.w(w127_19),.acc(r127_19),.res(r127_20),.clk(clk),.wout(w127_20));
	PE pe127_21(.x(x21),.w(w127_20),.acc(r127_20),.res(r127_21),.clk(clk),.wout(w127_21));
	PE pe127_22(.x(x22),.w(w127_21),.acc(r127_21),.res(r127_22),.clk(clk),.wout(w127_22));
	PE pe127_23(.x(x23),.w(w127_22),.acc(r127_22),.res(r127_23),.clk(clk),.wout(w127_23));
	PE pe127_24(.x(x24),.w(w127_23),.acc(r127_23),.res(r127_24),.clk(clk),.wout(w127_24));
	PE pe127_25(.x(x25),.w(w127_24),.acc(r127_24),.res(r127_25),.clk(clk),.wout(w127_25));
	PE pe127_26(.x(x26),.w(w127_25),.acc(r127_25),.res(r127_26),.clk(clk),.wout(w127_26));
	PE pe127_27(.x(x27),.w(w127_26),.acc(r127_26),.res(r127_27),.clk(clk),.wout(w127_27));
	PE pe127_28(.x(x28),.w(w127_27),.acc(r127_27),.res(r127_28),.clk(clk),.wout(w127_28));
	PE pe127_29(.x(x29),.w(w127_28),.acc(r127_28),.res(r127_29),.clk(clk),.wout(w127_29));
	PE pe127_30(.x(x30),.w(w127_29),.acc(r127_29),.res(r127_30),.clk(clk),.wout(w127_30));
	PE pe127_31(.x(x31),.w(w127_30),.acc(r127_30),.res(r127_31),.clk(clk),.wout(w127_31));
	PE pe127_32(.x(x32),.w(w127_31),.acc(r127_31),.res(r127_32),.clk(clk),.wout(w127_32));
	PE pe127_33(.x(x33),.w(w127_32),.acc(r127_32),.res(r127_33),.clk(clk),.wout(w127_33));
	PE pe127_34(.x(x34),.w(w127_33),.acc(r127_33),.res(r127_34),.clk(clk),.wout(w127_34));
	PE pe127_35(.x(x35),.w(w127_34),.acc(r127_34),.res(r127_35),.clk(clk),.wout(w127_35));
	PE pe127_36(.x(x36),.w(w127_35),.acc(r127_35),.res(r127_36),.clk(clk),.wout(w127_36));
	PE pe127_37(.x(x37),.w(w127_36),.acc(r127_36),.res(r127_37),.clk(clk),.wout(w127_37));
	PE pe127_38(.x(x38),.w(w127_37),.acc(r127_37),.res(r127_38),.clk(clk),.wout(w127_38));
	PE pe127_39(.x(x39),.w(w127_38),.acc(r127_38),.res(r127_39),.clk(clk),.wout(w127_39));
	PE pe127_40(.x(x40),.w(w127_39),.acc(r127_39),.res(r127_40),.clk(clk),.wout(w127_40));
	PE pe127_41(.x(x41),.w(w127_40),.acc(r127_40),.res(r127_41),.clk(clk),.wout(w127_41));
	PE pe127_42(.x(x42),.w(w127_41),.acc(r127_41),.res(r127_42),.clk(clk),.wout(w127_42));
	PE pe127_43(.x(x43),.w(w127_42),.acc(r127_42),.res(r127_43),.clk(clk),.wout(w127_43));
	PE pe127_44(.x(x44),.w(w127_43),.acc(r127_43),.res(r127_44),.clk(clk),.wout(w127_44));
	PE pe127_45(.x(x45),.w(w127_44),.acc(r127_44),.res(r127_45),.clk(clk),.wout(w127_45));
	PE pe127_46(.x(x46),.w(w127_45),.acc(r127_45),.res(r127_46),.clk(clk),.wout(w127_46));
	PE pe127_47(.x(x47),.w(w127_46),.acc(r127_46),.res(r127_47),.clk(clk),.wout(w127_47));
	PE pe127_48(.x(x48),.w(w127_47),.acc(r127_47),.res(r127_48),.clk(clk),.wout(w127_48));
	PE pe127_49(.x(x49),.w(w127_48),.acc(r127_48),.res(r127_49),.clk(clk),.wout(w127_49));
	PE pe127_50(.x(x50),.w(w127_49),.acc(r127_49),.res(r127_50),.clk(clk),.wout(w127_50));
	PE pe127_51(.x(x51),.w(w127_50),.acc(r127_50),.res(r127_51),.clk(clk),.wout(w127_51));
	PE pe127_52(.x(x52),.w(w127_51),.acc(r127_51),.res(r127_52),.clk(clk),.wout(w127_52));
	PE pe127_53(.x(x53),.w(w127_52),.acc(r127_52),.res(r127_53),.clk(clk),.wout(w127_53));
	PE pe127_54(.x(x54),.w(w127_53),.acc(r127_53),.res(r127_54),.clk(clk),.wout(w127_54));
	PE pe127_55(.x(x55),.w(w127_54),.acc(r127_54),.res(r127_55),.clk(clk),.wout(w127_55));
	PE pe127_56(.x(x56),.w(w127_55),.acc(r127_55),.res(r127_56),.clk(clk),.wout(w127_56));
	PE pe127_57(.x(x57),.w(w127_56),.acc(r127_56),.res(r127_57),.clk(clk),.wout(w127_57));
	PE pe127_58(.x(x58),.w(w127_57),.acc(r127_57),.res(r127_58),.clk(clk),.wout(w127_58));
	PE pe127_59(.x(x59),.w(w127_58),.acc(r127_58),.res(r127_59),.clk(clk),.wout(w127_59));
	PE pe127_60(.x(x60),.w(w127_59),.acc(r127_59),.res(r127_60),.clk(clk),.wout(w127_60));
	PE pe127_61(.x(x61),.w(w127_60),.acc(r127_60),.res(r127_61),.clk(clk),.wout(w127_61));
	PE pe127_62(.x(x62),.w(w127_61),.acc(r127_61),.res(r127_62),.clk(clk),.wout(w127_62));
	PE pe127_63(.x(x63),.w(w127_62),.acc(r127_62),.res(r127_63),.clk(clk),.wout(w127_63));
	PE pe127_64(.x(x64),.w(w127_63),.acc(r127_63),.res(r127_64),.clk(clk),.wout(w127_64));
	PE pe127_65(.x(x65),.w(w127_64),.acc(r127_64),.res(r127_65),.clk(clk),.wout(w127_65));
	PE pe127_66(.x(x66),.w(w127_65),.acc(r127_65),.res(r127_66),.clk(clk),.wout(w127_66));
	PE pe127_67(.x(x67),.w(w127_66),.acc(r127_66),.res(r127_67),.clk(clk),.wout(w127_67));
	PE pe127_68(.x(x68),.w(w127_67),.acc(r127_67),.res(r127_68),.clk(clk),.wout(w127_68));
	PE pe127_69(.x(x69),.w(w127_68),.acc(r127_68),.res(r127_69),.clk(clk),.wout(w127_69));
	PE pe127_70(.x(x70),.w(w127_69),.acc(r127_69),.res(r127_70),.clk(clk),.wout(w127_70));
	PE pe127_71(.x(x71),.w(w127_70),.acc(r127_70),.res(r127_71),.clk(clk),.wout(w127_71));
	PE pe127_72(.x(x72),.w(w127_71),.acc(r127_71),.res(r127_72),.clk(clk),.wout(w127_72));
	PE pe127_73(.x(x73),.w(w127_72),.acc(r127_72),.res(r127_73),.clk(clk),.wout(w127_73));
	PE pe127_74(.x(x74),.w(w127_73),.acc(r127_73),.res(r127_74),.clk(clk),.wout(w127_74));
	PE pe127_75(.x(x75),.w(w127_74),.acc(r127_74),.res(r127_75),.clk(clk),.wout(w127_75));
	PE pe127_76(.x(x76),.w(w127_75),.acc(r127_75),.res(r127_76),.clk(clk),.wout(w127_76));
	PE pe127_77(.x(x77),.w(w127_76),.acc(r127_76),.res(r127_77),.clk(clk),.wout(w127_77));
	PE pe127_78(.x(x78),.w(w127_77),.acc(r127_77),.res(r127_78),.clk(clk),.wout(w127_78));
	PE pe127_79(.x(x79),.w(w127_78),.acc(r127_78),.res(r127_79),.clk(clk),.wout(w127_79));
	PE pe127_80(.x(x80),.w(w127_79),.acc(r127_79),.res(r127_80),.clk(clk),.wout(w127_80));
	PE pe127_81(.x(x81),.w(w127_80),.acc(r127_80),.res(r127_81),.clk(clk),.wout(w127_81));
	PE pe127_82(.x(x82),.w(w127_81),.acc(r127_81),.res(r127_82),.clk(clk),.wout(w127_82));
	PE pe127_83(.x(x83),.w(w127_82),.acc(r127_82),.res(r127_83),.clk(clk),.wout(w127_83));
	PE pe127_84(.x(x84),.w(w127_83),.acc(r127_83),.res(r127_84),.clk(clk),.wout(w127_84));
	PE pe127_85(.x(x85),.w(w127_84),.acc(r127_84),.res(r127_85),.clk(clk),.wout(w127_85));
	PE pe127_86(.x(x86),.w(w127_85),.acc(r127_85),.res(r127_86),.clk(clk),.wout(w127_86));
	PE pe127_87(.x(x87),.w(w127_86),.acc(r127_86),.res(r127_87),.clk(clk),.wout(w127_87));
	PE pe127_88(.x(x88),.w(w127_87),.acc(r127_87),.res(r127_88),.clk(clk),.wout(w127_88));
	PE pe127_89(.x(x89),.w(w127_88),.acc(r127_88),.res(r127_89),.clk(clk),.wout(w127_89));
	PE pe127_90(.x(x90),.w(w127_89),.acc(r127_89),.res(r127_90),.clk(clk),.wout(w127_90));
	PE pe127_91(.x(x91),.w(w127_90),.acc(r127_90),.res(r127_91),.clk(clk),.wout(w127_91));
	PE pe127_92(.x(x92),.w(w127_91),.acc(r127_91),.res(r127_92),.clk(clk),.wout(w127_92));
	PE pe127_93(.x(x93),.w(w127_92),.acc(r127_92),.res(r127_93),.clk(clk),.wout(w127_93));
	PE pe127_94(.x(x94),.w(w127_93),.acc(r127_93),.res(r127_94),.clk(clk),.wout(w127_94));
	PE pe127_95(.x(x95),.w(w127_94),.acc(r127_94),.res(r127_95),.clk(clk),.wout(w127_95));
	PE pe127_96(.x(x96),.w(w127_95),.acc(r127_95),.res(r127_96),.clk(clk),.wout(w127_96));
	PE pe127_97(.x(x97),.w(w127_96),.acc(r127_96),.res(r127_97),.clk(clk),.wout(w127_97));
	PE pe127_98(.x(x98),.w(w127_97),.acc(r127_97),.res(r127_98),.clk(clk),.wout(w127_98));
	PE pe127_99(.x(x99),.w(w127_98),.acc(r127_98),.res(r127_99),.clk(clk),.wout(w127_99));
	PE pe127_100(.x(x100),.w(w127_99),.acc(r127_99),.res(r127_100),.clk(clk),.wout(w127_100));
	PE pe127_101(.x(x101),.w(w127_100),.acc(r127_100),.res(r127_101),.clk(clk),.wout(w127_101));
	PE pe127_102(.x(x102),.w(w127_101),.acc(r127_101),.res(r127_102),.clk(clk),.wout(w127_102));
	PE pe127_103(.x(x103),.w(w127_102),.acc(r127_102),.res(r127_103),.clk(clk),.wout(w127_103));
	PE pe127_104(.x(x104),.w(w127_103),.acc(r127_103),.res(r127_104),.clk(clk),.wout(w127_104));
	PE pe127_105(.x(x105),.w(w127_104),.acc(r127_104),.res(r127_105),.clk(clk),.wout(w127_105));
	PE pe127_106(.x(x106),.w(w127_105),.acc(r127_105),.res(r127_106),.clk(clk),.wout(w127_106));
	PE pe127_107(.x(x107),.w(w127_106),.acc(r127_106),.res(r127_107),.clk(clk),.wout(w127_107));
	PE pe127_108(.x(x108),.w(w127_107),.acc(r127_107),.res(r127_108),.clk(clk),.wout(w127_108));
	PE pe127_109(.x(x109),.w(w127_108),.acc(r127_108),.res(r127_109),.clk(clk),.wout(w127_109));
	PE pe127_110(.x(x110),.w(w127_109),.acc(r127_109),.res(r127_110),.clk(clk),.wout(w127_110));
	PE pe127_111(.x(x111),.w(w127_110),.acc(r127_110),.res(r127_111),.clk(clk),.wout(w127_111));
	PE pe127_112(.x(x112),.w(w127_111),.acc(r127_111),.res(r127_112),.clk(clk),.wout(w127_112));
	PE pe127_113(.x(x113),.w(w127_112),.acc(r127_112),.res(r127_113),.clk(clk),.wout(w127_113));
	PE pe127_114(.x(x114),.w(w127_113),.acc(r127_113),.res(r127_114),.clk(clk),.wout(w127_114));
	PE pe127_115(.x(x115),.w(w127_114),.acc(r127_114),.res(r127_115),.clk(clk),.wout(w127_115));
	PE pe127_116(.x(x116),.w(w127_115),.acc(r127_115),.res(r127_116),.clk(clk),.wout(w127_116));
	PE pe127_117(.x(x117),.w(w127_116),.acc(r127_116),.res(r127_117),.clk(clk),.wout(w127_117));
	PE pe127_118(.x(x118),.w(w127_117),.acc(r127_117),.res(r127_118),.clk(clk),.wout(w127_118));
	PE pe127_119(.x(x119),.w(w127_118),.acc(r127_118),.res(r127_119),.clk(clk),.wout(w127_119));
	PE pe127_120(.x(x120),.w(w127_119),.acc(r127_119),.res(r127_120),.clk(clk),.wout(w127_120));
	PE pe127_121(.x(x121),.w(w127_120),.acc(r127_120),.res(r127_121),.clk(clk),.wout(w127_121));
	PE pe127_122(.x(x122),.w(w127_121),.acc(r127_121),.res(r127_122),.clk(clk),.wout(w127_122));
	PE pe127_123(.x(x123),.w(w127_122),.acc(r127_122),.res(r127_123),.clk(clk),.wout(w127_123));
	PE pe127_124(.x(x124),.w(w127_123),.acc(r127_123),.res(r127_124),.clk(clk),.wout(w127_124));
	PE pe127_125(.x(x125),.w(w127_124),.acc(r127_124),.res(r127_125),.clk(clk),.wout(w127_125));
	PE pe127_126(.x(x126),.w(w127_125),.acc(r127_125),.res(r127_126),.clk(clk),.wout(w127_126));
	PE pe127_127(.x(x127),.w(w127_126),.acc(r127_126),.res(result127),.clk(clk),.wout(weight127));

endmodule